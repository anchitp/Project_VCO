* NGSPICE file created from Final_7_Flat.ext - technology: sky130A

.subckt Final_5_NSO VB OUT VP VCT VN
X0 a_6260_5590.t2 a_n1606_2236.t3 VP.t12 VP.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1 VP.t1 VCT.t0 a_9348_5588.t1 VP.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2 a_4518_1814.t1 a_1562_1830.t3 a_3194_252.t0 VN.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3 a_274_5606.t0 a_n1606_2236.t4 VP.t11 VP.t9 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4 a_4490_3828.t2 a_1534_3844.t3 a_9312_250.t1 VN.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5 a_3230_5590.t2 VCT.t1 VP.t4 VP.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6 a_n1698_2236.t1 a_n1698_2236.t0 VN.t11 VN.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=200000u
X7 a_n1606_2236.t1 a_n1606_2236.t0 VP.t10 VP.t9 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=200000u
X8 VP.t20 VCT.t2 a_12504_5562.t1 VP.t19 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9 a_12504_5562.t2 a_4518_1814.t3 OUT.t2 VP.t13 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10 a_6260_5590.t0 VCT.t3 VP.t3 VP.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X11 a_3230_5590.t0 a_4490_3828.t3 a_4518_1814.t2 VP.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X12 a_274_5606.t1 VCT.t4 VP.t14 VP.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X13 a_1562_1830.t1 a_1534_3844.t4 a_274_5606.t2 VP.t17 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X14 a_9312_250.t2 a_1976_242.t2 VN.t17 VN.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X15 a_12504_5562.t0 a_n1606_2236.t5 VP.t8 VP.t7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X16 a_1562_1830.t0 OUT.t3 a_238_268.t0 VN.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X17 a_12468_224.t1 a_1976_242.t3 VN.t19 VN.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X18 a_9348_5588.t0 a_n1606_2236.t6 VP.t6 VP.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X19 a_1534_3844.t1 OUT.t4 a_6260_5590.t1 VP.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X20 VN.t5 a_n1698_2236.t3 a_6224_252.t1 VN.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X21 a_n1698_2236.t2 VB.t0 a_n1606_2236.t2 VN.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X22 a_1534_3844.t2 a_4518_1814.t4 a_6224_252.t2 VN.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X23 a_6224_252.t0 a_1976_242.t4 VN.t18 VN.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X24 a_3230_5590.t1 a_n1606_2236.t7 VP.t5 VP.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X25 a_3194_252.t2 a_1976_242.t5 VN.t21 VN.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X26 OUT.t0 a_4490_3828.t4 a_12468_224.t0 VN.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X27 a_9312_250.t0 a_n1698_2236.t4 VN.t6 VN.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X28 a_9348_5588.t2 a_1562_1830.t4 a_4490_3828.t0 VP.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X29 VN.t7 a_n1698_2236.t5 a_12468_224.t2 VN.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X30 a_1534_3844.t0 OUT.t5 VN.t10 VN.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X31 VN.t22 a_1976_242.t6 a_238_268.t1 VN.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X32 VN.t12 a_n1698_2236.t6 a_3194_252.t1 VN.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X33 OUT.t1 a_4518_1814.t5 VN.t15 VN.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X34 a_4518_1814.t0 a_4490_3828.t5 VN.t3 VN.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X35 a_238_268.t2 a_n1698_2236.t7 VN.t13 VN.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X36 VP.t16 VN.t23 a_1976_242.t1 VP.t15 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X37 a_1976_242.t0 VCT.t5 VN.t14 VN.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X38 a_4490_3828.t1 a_1562_1830.t5 VN.t8 VN.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X39 a_1562_1830.t2 a_1534_3844.t5 VN.t16 VN.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
R0 a_n1606_2236.n50 a_n1606_2236.n49 1018.63
R1 a_n1606_2236.n72 a_n1606_2236.n71 1018.63
R2 a_n1606_2236.n94 a_n1606_2236.n93 1018.63
R3 a_n1606_2236.n116 a_n1606_2236.n115 1018.63
R4 a_n1606_2236.n138 a_n1606_2236.n137 1018.63
R5 a_n1606_2236.n61 a_n1606_2236.n60 926.657
R6 a_n1606_2236.n83 a_n1606_2236.n82 926.657
R7 a_n1606_2236.n105 a_n1606_2236.n104 926.657
R8 a_n1606_2236.n127 a_n1606_2236.n126 926.657
R9 a_n1606_2236.n149 a_n1606_2236.n148 926.657
R10 a_n1606_2236.n58 a_n1606_2236.t4 864.386
R11 a_n1606_2236.n57 a_n1606_2236.n41 864.386
R12 a_n1606_2236.n56 a_n1606_2236.n42 864.386
R13 a_n1606_2236.n55 a_n1606_2236.n43 864.386
R14 a_n1606_2236.n54 a_n1606_2236.n44 864.386
R15 a_n1606_2236.n53 a_n1606_2236.n45 864.386
R16 a_n1606_2236.n52 a_n1606_2236.n46 864.386
R17 a_n1606_2236.n51 a_n1606_2236.n47 864.386
R18 a_n1606_2236.n50 a_n1606_2236.n48 864.386
R19 a_n1606_2236.n59 a_n1606_2236.n40 864.386
R20 a_n1606_2236.n80 a_n1606_2236.n63 864.386
R21 a_n1606_2236.n79 a_n1606_2236.n64 864.386
R22 a_n1606_2236.n78 a_n1606_2236.n65 864.386
R23 a_n1606_2236.n77 a_n1606_2236.n66 864.386
R24 a_n1606_2236.n76 a_n1606_2236.n67 864.386
R25 a_n1606_2236.n75 a_n1606_2236.n68 864.386
R26 a_n1606_2236.n74 a_n1606_2236.n69 864.386
R27 a_n1606_2236.n73 a_n1606_2236.n70 864.386
R28 a_n1606_2236.n72 a_n1606_2236.t7 864.386
R29 a_n1606_2236.n81 a_n1606_2236.n62 864.386
R30 a_n1606_2236.n102 a_n1606_2236.n85 864.386
R31 a_n1606_2236.n101 a_n1606_2236.n86 864.386
R32 a_n1606_2236.n100 a_n1606_2236.n87 864.386
R33 a_n1606_2236.n99 a_n1606_2236.n88 864.386
R34 a_n1606_2236.n98 a_n1606_2236.n89 864.386
R35 a_n1606_2236.n97 a_n1606_2236.n90 864.386
R36 a_n1606_2236.n96 a_n1606_2236.n91 864.386
R37 a_n1606_2236.n95 a_n1606_2236.n92 864.386
R38 a_n1606_2236.n94 a_n1606_2236.t3 864.386
R39 a_n1606_2236.n103 a_n1606_2236.n84 864.386
R40 a_n1606_2236.n124 a_n1606_2236.n107 864.386
R41 a_n1606_2236.n123 a_n1606_2236.n108 864.386
R42 a_n1606_2236.n122 a_n1606_2236.n109 864.386
R43 a_n1606_2236.n121 a_n1606_2236.n110 864.386
R44 a_n1606_2236.n120 a_n1606_2236.t6 864.386
R45 a_n1606_2236.n119 a_n1606_2236.n111 864.386
R46 a_n1606_2236.n118 a_n1606_2236.n112 864.386
R47 a_n1606_2236.n117 a_n1606_2236.n113 864.386
R48 a_n1606_2236.n116 a_n1606_2236.n114 864.386
R49 a_n1606_2236.n125 a_n1606_2236.n106 864.386
R50 a_n1606_2236.n146 a_n1606_2236.t5 864.386
R51 a_n1606_2236.n145 a_n1606_2236.n129 864.386
R52 a_n1606_2236.n144 a_n1606_2236.n130 864.386
R53 a_n1606_2236.n143 a_n1606_2236.n131 864.386
R54 a_n1606_2236.n142 a_n1606_2236.n132 864.386
R55 a_n1606_2236.n141 a_n1606_2236.n133 864.386
R56 a_n1606_2236.n140 a_n1606_2236.n134 864.386
R57 a_n1606_2236.n139 a_n1606_2236.n135 864.386
R58 a_n1606_2236.n138 a_n1606_2236.n136 864.386
R59 a_n1606_2236.n147 a_n1606_2236.n128 864.386
R60 a_n1606_2236.n166 a_n1606_2236.n165 783.313
R61 a_n1606_2236.n157 a_n1606_2236.n155 783.313
R62 a_n1606_2236.n166 a_n1606_2236.t0 709.745
R63 a_n1606_2236.n157 a_n1606_2236.n156 709.745
R64 a_n1606_2236.n160 a_n1606_2236.n159 709.745
R65 a_n1606_2236.n162 a_n1606_2236.n161 709.745
R66 a_n1606_2236.n164 a_n1606_2236.n163 709.745
R67 a_n1606_2236.n158 a_n1606_2236.n154 684.44
R68 a_n1606_2236.n193 a_n1606_2236.n183 281.697
R69 a_n1606_2236.n150 a_n1606_2236.n149 204.487
R70 a_n1606_2236.n150 a_n1606_2236.n127 202.574
R71 a_n1606_2236.n152 a_n1606_2236.n83 202.57
R72 a_n1606_2236.n151 a_n1606_2236.n105 202.57
R73 a_n1606_2236.n153 a_n1606_2236.n61 202.538
R74 a_n1606_2236.n51 a_n1606_2236.n50 154.24
R75 a_n1606_2236.n52 a_n1606_2236.n51 154.24
R76 a_n1606_2236.n53 a_n1606_2236.n52 154.24
R77 a_n1606_2236.n54 a_n1606_2236.n53 154.24
R78 a_n1606_2236.n55 a_n1606_2236.n54 154.24
R79 a_n1606_2236.n56 a_n1606_2236.n55 154.24
R80 a_n1606_2236.n57 a_n1606_2236.n56 154.24
R81 a_n1606_2236.n58 a_n1606_2236.n57 154.24
R82 a_n1606_2236.n73 a_n1606_2236.n72 154.24
R83 a_n1606_2236.n74 a_n1606_2236.n73 154.24
R84 a_n1606_2236.n75 a_n1606_2236.n74 154.24
R85 a_n1606_2236.n76 a_n1606_2236.n75 154.24
R86 a_n1606_2236.n77 a_n1606_2236.n76 154.24
R87 a_n1606_2236.n78 a_n1606_2236.n77 154.24
R88 a_n1606_2236.n79 a_n1606_2236.n78 154.24
R89 a_n1606_2236.n80 a_n1606_2236.n79 154.24
R90 a_n1606_2236.n95 a_n1606_2236.n94 154.24
R91 a_n1606_2236.n96 a_n1606_2236.n95 154.24
R92 a_n1606_2236.n97 a_n1606_2236.n96 154.24
R93 a_n1606_2236.n98 a_n1606_2236.n97 154.24
R94 a_n1606_2236.n99 a_n1606_2236.n98 154.24
R95 a_n1606_2236.n100 a_n1606_2236.n99 154.24
R96 a_n1606_2236.n101 a_n1606_2236.n100 154.24
R97 a_n1606_2236.n102 a_n1606_2236.n101 154.24
R98 a_n1606_2236.n117 a_n1606_2236.n116 154.24
R99 a_n1606_2236.n118 a_n1606_2236.n117 154.24
R100 a_n1606_2236.n119 a_n1606_2236.n118 154.24
R101 a_n1606_2236.n120 a_n1606_2236.n119 154.24
R102 a_n1606_2236.n121 a_n1606_2236.n120 154.24
R103 a_n1606_2236.n122 a_n1606_2236.n121 154.24
R104 a_n1606_2236.n123 a_n1606_2236.n122 154.24
R105 a_n1606_2236.n124 a_n1606_2236.n123 154.24
R106 a_n1606_2236.n139 a_n1606_2236.n138 154.24
R107 a_n1606_2236.n140 a_n1606_2236.n139 154.24
R108 a_n1606_2236.n141 a_n1606_2236.n140 154.24
R109 a_n1606_2236.n142 a_n1606_2236.n141 154.24
R110 a_n1606_2236.n143 a_n1606_2236.n142 154.24
R111 a_n1606_2236.n144 a_n1606_2236.n143 154.24
R112 a_n1606_2236.n145 a_n1606_2236.n144 154.24
R113 a_n1606_2236.n146 a_n1606_2236.n145 154.24
R114 a_n1606_2236.n59 a_n1606_2236.n58 142.605
R115 a_n1606_2236.n81 a_n1606_2236.n80 142.605
R116 a_n1606_2236.n103 a_n1606_2236.n102 142.605
R117 a_n1606_2236.n125 a_n1606_2236.n124 142.605
R118 a_n1606_2236.n147 a_n1606_2236.n146 142.605
R119 a_n1606_2236.n179 a_n1606_2236.n178 115.46
R120 a_n1606_2236.n181 a_n1606_2236.n169 113.686
R121 a_n1606_2236.n182 a_n1606_2236.n167 112.463
R122 a_n1606_2236.n160 a_n1606_2236.n158 97.668
R123 a_n1606_2236.n158 a_n1606_2236.n157 97.541
R124 a_n1606_2236.n183 a_n1606_2236.n182 76
R125 a_n1606_2236.n162 a_n1606_2236.n160 73.568
R126 a_n1606_2236.n164 a_n1606_2236.n162 73.568
R127 a_n1606_2236.n180 a_n1606_2236.n179 69.99
R128 a_n1606_2236.n182 a_n1606_2236.n181 58.332
R129 a_n1606_2236.t2 a_n1606_2236.n193 122.225
R130 a_n1606_2236.n179 a_n1606_2236.n175 45.131
R131 a_n1606_2236.n180 a_n1606_2236.n172 45.131
R132 a_n1606_2236.n61 a_n1606_2236.n59 41.551
R133 a_n1606_2236.n83 a_n1606_2236.n81 41.551
R134 a_n1606_2236.n105 a_n1606_2236.n103 41.551
R135 a_n1606_2236.n127 a_n1606_2236.n125 41.551
R136 a_n1606_2236.n149 a_n1606_2236.n147 41.551
R137 a_n1606_2236.t2 a_n1606_2236.n39 32.727
R138 a_n1606_2236.n39 a_n1606_2236.n1 29.09
R139 a_n1606_2236.n187 a_n1606_2236.n186 20
R140 a_n1606_2236.n6 a_n1606_2236.n5 16.363
R141 a_n1606_2236.n167 a_n1606_2236.n166 15.221
R142 a_n1606_2236.n31 a_n1606_2236.n30 15
R143 a_n1606_2236.n23 a_n1606_2236.n22 15
R144 a_n1606_2236.n15 a_n1606_2236.n14 15
R145 a_n1606_2236.n7 a_n1606_2236.n6 15
R146 a_n1606_2236.n188 a_n1606_2236.n187 15
R147 a_n1606_2236.n39 a_n1606_2236.n38 15
R148 a_n1606_2236.n33 a_n1606_2236.n32 15
R149 a_n1606_2236.n25 a_n1606_2236.n24 15
R150 a_n1606_2236.n17 a_n1606_2236.n16 15
R151 a_n1606_2236.n9 a_n1606_2236.n8 15
R152 a_n1606_2236.n185 a_n1606_2236.n184 15
R153 a_n1606_2236.n192 a_n1606_2236.n191 13.634
R154 a_n1606_2236.n10 a_n1606_2236.n9 12.917
R155 a_n1606_2236.n18 a_n1606_2236.n17 12.917
R156 a_n1606_2236.n26 a_n1606_2236.n25 12.917
R157 a_n1606_2236.n34 a_n1606_2236.n33 12.917
R158 a_n1606_2236.n14 a_n1606_2236.n13 12.727
R159 a_n1606_2236.n22 a_n1606_2236.n21 9.09
R160 a_n1606_2236.n193 a_n1606_2236.n192 8.695
R161 a_n1606_2236.n167 a_n1606_2236.n164 7.61
R162 a_n1606_2236.n35 a_n1606_2236.n34 5.741
R163 a_n1606_2236.n38 a_n1606_2236.n37 5.741
R164 a_n1606_2236.n175 a_n1606_2236.n173 5.713
R165 a_n1606_2236.n175 a_n1606_2236.n174 5.713
R166 a_n1606_2236.n178 a_n1606_2236.n176 5.713
R167 a_n1606_2236.n178 a_n1606_2236.n177 5.713
R168 a_n1606_2236.n169 a_n1606_2236.n168 5.713
R169 a_n1606_2236.n169 a_n1606_2236.t1 5.713
R170 a_n1606_2236.n172 a_n1606_2236.n170 5.713
R171 a_n1606_2236.n172 a_n1606_2236.n171 5.713
R172 a_n1606_2236.n30 a_n1606_2236.n29 5.454
R173 a_n1606_2236.n27 a_n1606_2236.n26 5.023
R174 a_n1606_2236.n33 a_n1606_2236.n31 5.023
R175 a_n1606_2236.n19 a_n1606_2236.n18 4.305
R176 a_n1606_2236.n25 a_n1606_2236.n23 4.305
R177 a_n1606_2236.n190 a_n1606_2236.n189 3.947
R178 a_n1606_2236.n189 a_n1606_2236.n188 3.947
R179 a_n1606_2236.n11 a_n1606_2236.n10 3.588
R180 a_n1606_2236.n17 a_n1606_2236.n15 3.588
R181 a_n1606_2236.n4 a_n1606_2236.n3 3.229
R182 a_n1606_2236.n7 a_n1606_2236.n4 3.229
R183 a_n1606_2236.n3 a_n1606_2236.n2 2.87
R184 a_n1606_2236.n9 a_n1606_2236.n7 2.87
R185 a_n1606_2236.n183 a_n1606_2236.n153 2.668
R186 a_n1606_2236.n12 a_n1606_2236.n11 2.511
R187 a_n1606_2236.n15 a_n1606_2236.n12 2.511
R188 a_n1606_2236.n191 a_n1606_2236.n190 2.152
R189 a_n1606_2236.n188 a_n1606_2236.n185 2.152
R190 a_n1606_2236.n151 a_n1606_2236.n150 1.82
R191 a_n1606_2236.n1 a_n1606_2236.n0 1.818
R192 a_n1606_2236.n20 a_n1606_2236.n19 1.794
R193 a_n1606_2236.n23 a_n1606_2236.n20 1.794
R194 a_n1606_2236.n152 a_n1606_2236.n151 1.786
R195 a_n1606_2236.n153 a_n1606_2236.n152 1.742
R196 a_n1606_2236.n181 a_n1606_2236.n180 1.355
R197 a_n1606_2236.n28 a_n1606_2236.n27 1.076
R198 a_n1606_2236.n31 a_n1606_2236.n28 1.076
R199 a_n1606_2236.n36 a_n1606_2236.n35 0.358
R200 a_n1606_2236.n37 a_n1606_2236.n36 0.358
R201 VP.n766 VP.t9 530.876
R202 VP.t7 VP.t13 442.607
R203 VP.t0 VP.t7 408.504
R204 VP.t13 VP.t19 389.969
R205 VP.t2 VP.t18 371.434
R206 VP.n558 VP.n557 314.834
R207 VP.n138 VP.n137 314.754
R208 VP.n558 VP.n488 310.804
R209 VP.n416 VP.n415 310.491
R210 VP.t17 VP.t2 289.379
R211 VP.t19 VP.t15 278.761
R212 VP.t18 VP.t0 247.623
R213 VP.n416 VP.n346 241.911
R214 VP.n767 VP.n766 218.582
R215 VP.n417 VP.t16 212.355
R216 VP.n768 VP.n767 185.797
R217 VP.n277 VP.n276 176.93
R218 VP.n277 VP.n207 173.108
R219 VP.n138 VP.n68 173.066
R220 VP.n768 VP.n627 172.942
R221 VP.n766 VP.n765 150.175
R222 VP.n712 VP.t10 72.48
R223 VP.n435 VP.t4 68.375
R224 VP.n293 VP.t20 68.375
R225 VP.n643 VP.t11 64.755
R226 VP.n574 VP.t14 64.755
R227 VP.n504 VP.t5 64.755
R228 VP.n84 VP.t12 64.755
R229 VP.n15 VP.t3 64.755
R230 VP.n223 VP.t6 64.755
R231 VP.n154 VP.t1 64.755
R232 VP.n362 VP.t8 64.755
R233 VP.n765 VP.n730 49.503
R234 VP.n696 VP.n661 49.503
R235 VP.n627 VP.n592 49.503
R236 VP.n557 VP.n522 49.503
R237 VP.n488 VP.n453 49.503
R238 VP.n137 VP.n102 49.503
R239 VP.n68 VP.n33 49.503
R240 VP.n276 VP.n241 49.503
R241 VP.n207 VP.n172 49.503
R242 VP.n415 VP.n380 49.503
R243 VP.n346 VP.n311 49.503
R244 VP.n759 VP.n758 37.362
R245 VP.n482 VP.n481 34.951
R246 VP.n340 VP.n339 34.951
R247 VP.n690 VP.n689 32.833
R248 VP.n621 VP.n620 32.833
R249 VP.n551 VP.n550 32.833
R250 VP.n131 VP.n130 32.833
R251 VP.n62 VP.n61 32.833
R252 VP.n270 VP.n269 32.833
R253 VP.n201 VP.n200 32.833
R254 VP.n409 VP.n408 32.833
R255 VP.n713 VP.n712 30.824
R256 VP.n436 VP.n435 30.687
R257 VP.n294 VP.n293 30.687
R258 VP.n751 VP.n750 30.568
R259 VP.n644 VP.n643 30.553
R260 VP.n575 VP.n574 30.553
R261 VP.n505 VP.n504 30.553
R262 VP.n85 VP.n84 30.553
R263 VP.n16 VP.n15 30.553
R264 VP.n224 VP.n223 30.553
R265 VP.n155 VP.n154 30.553
R266 VP.n363 VP.n362 30.553
R267 VP.n474 VP.n473 28.596
R268 VP.n332 VP.n331 28.596
R269 VP.n682 VP.n681 26.863
R270 VP.n613 VP.n612 26.863
R271 VP.n543 VP.n542 26.863
R272 VP.n123 VP.n122 26.863
R273 VP.n54 VP.n53 26.863
R274 VP.n262 VP.n261 26.863
R275 VP.n193 VP.n192 26.863
R276 VP.n401 VP.n400 26.863
R277 VP.n767 VP.n696 26.144
R278 VP.n743 VP.n742 23.775
R279 VP.n466 VP.n465 22.241
R280 VP.n324 VP.n323 22.241
R281 VP.n674 VP.n673 20.893
R282 VP.n605 VP.n604 20.893
R283 VP.n535 VP.n534 20.893
R284 VP.n115 VP.n114 20.893
R285 VP.n46 VP.n45 20.893
R286 VP.n254 VP.n253 20.893
R287 VP.n185 VP.n184 20.893
R288 VP.n393 VP.n392 20.893
R289 VP.n735 VP.n734 16.982
R290 VP.n458 VP.n457 15.887
R291 VP.n316 VP.n315 15.887
R292 VP.n709 VP.n708 15
R293 VP.n701 VP.n700 15
R294 VP.n736 VP.n735 15
R295 VP.n744 VP.n743 15
R296 VP.n752 VP.n751 15
R297 VP.n760 VP.n759 15
R298 VP.n711 VP.n710 15
R299 VP.n703 VP.n702 15
R300 VP.n733 VP.n732 15
R301 VP.n741 VP.n740 15
R302 VP.n749 VP.n748 15
R303 VP.n757 VP.n756 15
R304 VP.n640 VP.n639 15
R305 VP.n632 VP.n631 15
R306 VP.n667 VP.n666 15
R307 VP.n675 VP.n674 15
R308 VP.n683 VP.n682 15
R309 VP.n691 VP.n690 15
R310 VP.n642 VP.n641 15
R311 VP.n634 VP.n633 15
R312 VP.n664 VP.n663 15
R313 VP.n672 VP.n671 15
R314 VP.n680 VP.n679 15
R315 VP.n688 VP.n687 15
R316 VP.n571 VP.n570 15
R317 VP.n563 VP.n562 15
R318 VP.n598 VP.n597 15
R319 VP.n606 VP.n605 15
R320 VP.n614 VP.n613 15
R321 VP.n622 VP.n621 15
R322 VP.n573 VP.n572 15
R323 VP.n565 VP.n564 15
R324 VP.n595 VP.n594 15
R325 VP.n603 VP.n602 15
R326 VP.n611 VP.n610 15
R327 VP.n619 VP.n618 15
R328 VP.n501 VP.n500 15
R329 VP.n493 VP.n492 15
R330 VP.n528 VP.n527 15
R331 VP.n536 VP.n535 15
R332 VP.n544 VP.n543 15
R333 VP.n552 VP.n551 15
R334 VP.n503 VP.n502 15
R335 VP.n495 VP.n494 15
R336 VP.n525 VP.n524 15
R337 VP.n533 VP.n532 15
R338 VP.n541 VP.n540 15
R339 VP.n549 VP.n548 15
R340 VP.n432 VP.n431 15
R341 VP.n424 VP.n423 15
R342 VP.n459 VP.n458 15
R343 VP.n467 VP.n466 15
R344 VP.n475 VP.n474 15
R345 VP.n483 VP.n482 15
R346 VP.n434 VP.n433 15
R347 VP.n426 VP.n425 15
R348 VP.n456 VP.n455 15
R349 VP.n464 VP.n463 15
R350 VP.n472 VP.n471 15
R351 VP.n480 VP.n479 15
R352 VP.n81 VP.n80 15
R353 VP.n73 VP.n72 15
R354 VP.n108 VP.n107 15
R355 VP.n116 VP.n115 15
R356 VP.n124 VP.n123 15
R357 VP.n132 VP.n131 15
R358 VP.n83 VP.n82 15
R359 VP.n75 VP.n74 15
R360 VP.n105 VP.n104 15
R361 VP.n113 VP.n112 15
R362 VP.n121 VP.n120 15
R363 VP.n129 VP.n128 15
R364 VP.n12 VP.n11 15
R365 VP.n4 VP.n3 15
R366 VP.n39 VP.n38 15
R367 VP.n47 VP.n46 15
R368 VP.n55 VP.n54 15
R369 VP.n63 VP.n62 15
R370 VP.n14 VP.n13 15
R371 VP.n6 VP.n5 15
R372 VP.n36 VP.n35 15
R373 VP.n44 VP.n43 15
R374 VP.n52 VP.n51 15
R375 VP.n60 VP.n59 15
R376 VP.n220 VP.n219 15
R377 VP.n212 VP.n211 15
R378 VP.n247 VP.n246 15
R379 VP.n255 VP.n254 15
R380 VP.n263 VP.n262 15
R381 VP.n271 VP.n270 15
R382 VP.n222 VP.n221 15
R383 VP.n214 VP.n213 15
R384 VP.n244 VP.n243 15
R385 VP.n252 VP.n251 15
R386 VP.n260 VP.n259 15
R387 VP.n268 VP.n267 15
R388 VP.n151 VP.n150 15
R389 VP.n143 VP.n142 15
R390 VP.n178 VP.n177 15
R391 VP.n186 VP.n185 15
R392 VP.n194 VP.n193 15
R393 VP.n202 VP.n201 15
R394 VP.n153 VP.n152 15
R395 VP.n145 VP.n144 15
R396 VP.n175 VP.n174 15
R397 VP.n183 VP.n182 15
R398 VP.n191 VP.n190 15
R399 VP.n199 VP.n198 15
R400 VP.n359 VP.n358 15
R401 VP.n351 VP.n350 15
R402 VP.n386 VP.n385 15
R403 VP.n394 VP.n393 15
R404 VP.n402 VP.n401 15
R405 VP.n410 VP.n409 15
R406 VP.n361 VP.n360 15
R407 VP.n353 VP.n352 15
R408 VP.n383 VP.n382 15
R409 VP.n391 VP.n390 15
R410 VP.n399 VP.n398 15
R411 VP.n407 VP.n406 15
R412 VP.n290 VP.n289 15
R413 VP.n282 VP.n281 15
R414 VP.n317 VP.n316 15
R415 VP.n325 VP.n324 15
R416 VP.n333 VP.n332 15
R417 VP.n341 VP.n340 15
R418 VP.n292 VP.n291 15
R419 VP.n284 VP.n283 15
R420 VP.n314 VP.n313 15
R421 VP.n322 VP.n321 15
R422 VP.n330 VP.n329 15
R423 VP.n338 VP.n337 15
R424 VP.n666 VP.n665 14.924
R425 VP.n597 VP.n596 14.924
R426 VP.n527 VP.n526 14.924
R427 VP.n107 VP.n106 14.924
R428 VP.n38 VP.n37 14.924
R429 VP.n246 VP.n245 14.924
R430 VP.n177 VP.n176 14.924
R431 VP.n385 VP.n384 14.924
R432 VP.n643 VP.n642 14.123
R433 VP.n574 VP.n573 14.123
R434 VP.n504 VP.n503 14.123
R435 VP.n84 VP.n83 14.123
R436 VP.n15 VP.n14 14.123
R437 VP.n223 VP.n222 14.123
R438 VP.n154 VP.n153 14.123
R439 VP.n362 VP.n361 14.123
R440 VP.n435 VP.n434 14.071
R441 VP.n293 VP.n292 14.071
R442 VP.n712 VP.n711 14.017
R443 VP.n695 VP.n694 13.544
R444 VP.n626 VP.n625 13.544
R445 VP.n556 VP.n555 13.544
R446 VP.n136 VP.n135 13.544
R447 VP.n67 VP.n66 13.544
R448 VP.n275 VP.n274 13.544
R449 VP.n206 VP.n205 13.544
R450 VP.n414 VP.n413 13.544
R451 VP.n487 VP.n486 13.532
R452 VP.n345 VP.n344 13.532
R453 VP.n764 VP.n763 13.518
R454 VP.n757 VP.n755 12.917
R455 VP.n749 VP.n747 12.917
R456 VP.n741 VP.n739 12.917
R457 VP.n733 VP.n731 12.917
R458 VP.n704 VP.n703 12.917
R459 VP.n688 VP.n686 12.917
R460 VP.n680 VP.n678 12.917
R461 VP.n672 VP.n670 12.917
R462 VP.n664 VP.n662 12.917
R463 VP.n635 VP.n634 12.917
R464 VP.n619 VP.n617 12.917
R465 VP.n611 VP.n609 12.917
R466 VP.n603 VP.n601 12.917
R467 VP.n595 VP.n593 12.917
R468 VP.n566 VP.n565 12.917
R469 VP.n549 VP.n547 12.917
R470 VP.n541 VP.n539 12.917
R471 VP.n533 VP.n531 12.917
R472 VP.n525 VP.n523 12.917
R473 VP.n496 VP.n495 12.917
R474 VP.n480 VP.n478 12.917
R475 VP.n472 VP.n470 12.917
R476 VP.n464 VP.n462 12.917
R477 VP.n456 VP.n454 12.917
R478 VP.n427 VP.n426 12.917
R479 VP.n129 VP.n127 12.917
R480 VP.n121 VP.n119 12.917
R481 VP.n113 VP.n111 12.917
R482 VP.n105 VP.n103 12.917
R483 VP.n76 VP.n75 12.917
R484 VP.n60 VP.n58 12.917
R485 VP.n52 VP.n50 12.917
R486 VP.n44 VP.n42 12.917
R487 VP.n36 VP.n34 12.917
R488 VP.n7 VP.n6 12.917
R489 VP.n268 VP.n266 12.917
R490 VP.n260 VP.n258 12.917
R491 VP.n252 VP.n250 12.917
R492 VP.n244 VP.n242 12.917
R493 VP.n215 VP.n214 12.917
R494 VP.n199 VP.n197 12.917
R495 VP.n191 VP.n189 12.917
R496 VP.n183 VP.n181 12.917
R497 VP.n175 VP.n173 12.917
R498 VP.n146 VP.n145 12.917
R499 VP.n407 VP.n405 12.917
R500 VP.n399 VP.n397 12.917
R501 VP.n391 VP.n389 12.917
R502 VP.n383 VP.n381 12.917
R503 VP.n354 VP.n353 12.917
R504 VP.n338 VP.n336 12.917
R505 VP.n330 VP.n328 12.917
R506 VP.n322 VP.n320 12.917
R507 VP.n314 VP.n312 12.917
R508 VP.n285 VP.n284 12.917
R509 VP.n700 VP.n699 10.189
R510 VP.n423 VP.n422 9.532
R511 VP.n281 VP.n280 9.532
R512 VP.n631 VP.n630 8.954
R513 VP.n562 VP.n561 8.954
R514 VP.n492 VP.n491 8.954
R515 VP.n72 VP.n71 8.954
R516 VP.n3 VP.n2 8.954
R517 VP.n211 VP.n210 8.954
R518 VP.n142 VP.n141 8.954
R519 VP.n350 VP.n349 8.954
R520 VP.n765 VP.n764 8.838
R521 VP.n488 VP.n487 8.82
R522 VP.n346 VP.n345 8.82
R523 VP.n696 VP.n695 8.805
R524 VP.n627 VP.n626 8.805
R525 VP.n557 VP.n556 8.805
R526 VP.n137 VP.n136 8.805
R527 VP.n68 VP.n67 8.805
R528 VP.n276 VP.n275 8.805
R529 VP.n207 VP.n206 8.805
R530 VP.n415 VP.n414 8.805
R531 VP.t9 VP.t17 7.617
R532 VP.n769 VP.n558 6.506
R533 VP.n418 VP.n277 6.475
R534 VP.n419 VP.n138 6.473
R535 VP.n417 VP.n416 6.417
R536 VP.n705 VP.n704 5.741
R537 VP.n711 VP.n709 5.741
R538 VP.n636 VP.n635 5.741
R539 VP.n642 VP.n640 5.741
R540 VP.n567 VP.n566 5.741
R541 VP.n573 VP.n571 5.741
R542 VP.n497 VP.n496 5.741
R543 VP.n503 VP.n501 5.741
R544 VP.n428 VP.n427 5.741
R545 VP.n434 VP.n432 5.741
R546 VP.n77 VP.n76 5.741
R547 VP.n83 VP.n81 5.741
R548 VP.n8 VP.n7 5.741
R549 VP.n14 VP.n12 5.741
R550 VP.n216 VP.n215 5.741
R551 VP.n222 VP.n220 5.741
R552 VP.n147 VP.n146 5.741
R553 VP.n153 VP.n151 5.741
R554 VP.n355 VP.n354 5.741
R555 VP.n361 VP.n359 5.741
R556 VP.n286 VP.n285 5.741
R557 VP.n292 VP.n290 5.741
R558 VP.n703 VP.n701 5.023
R559 VP.n634 VP.n632 5.023
R560 VP.n565 VP.n563 5.023
R561 VP.n495 VP.n493 5.023
R562 VP.n426 VP.n424 5.023
R563 VP.n75 VP.n73 5.023
R564 VP.n6 VP.n4 5.023
R565 VP.n214 VP.n212 5.023
R566 VP.n145 VP.n143 5.023
R567 VP.n353 VP.n351 5.023
R568 VP.n284 VP.n282 5.023
R569 VP.n769 VP.n768 4.734
R570 VP.n739 VP.n738 4.305
R571 VP.n736 VP.n733 4.305
R572 VP.n670 VP.n669 4.305
R573 VP.n667 VP.n664 4.305
R574 VP.n601 VP.n600 4.305
R575 VP.n598 VP.n595 4.305
R576 VP.n531 VP.n530 4.305
R577 VP.n528 VP.n525 4.305
R578 VP.n462 VP.n461 4.305
R579 VP.n459 VP.n456 4.305
R580 VP.n111 VP.n110 4.305
R581 VP.n108 VP.n105 4.305
R582 VP.n42 VP.n41 4.305
R583 VP.n39 VP.n36 4.305
R584 VP.n250 VP.n249 4.305
R585 VP.n247 VP.n244 4.305
R586 VP.n181 VP.n180 4.305
R587 VP.n178 VP.n175 4.305
R588 VP.n389 VP.n388 4.305
R589 VP.n386 VP.n383 4.305
R590 VP.n320 VP.n319 4.305
R591 VP.n317 VP.n314 4.305
R592 VP.n762 VP.n761 3.947
R593 VP.n761 VP.n760 3.947
R594 VP.n693 VP.n692 3.947
R595 VP.n692 VP.n691 3.947
R596 VP.n624 VP.n623 3.947
R597 VP.n623 VP.n622 3.947
R598 VP.n554 VP.n553 3.947
R599 VP.n553 VP.n552 3.947
R600 VP.n485 VP.n484 3.947
R601 VP.n484 VP.n483 3.947
R602 VP.n134 VP.n133 3.947
R603 VP.n133 VP.n132 3.947
R604 VP.n65 VP.n64 3.947
R605 VP.n64 VP.n63 3.947
R606 VP.n273 VP.n272 3.947
R607 VP.n272 VP.n271 3.947
R608 VP.n204 VP.n203 3.947
R609 VP.n203 VP.n202 3.947
R610 VP.n412 VP.n411 3.947
R611 VP.n411 VP.n410 3.947
R612 VP.n343 VP.n342 3.947
R613 VP.n342 VP.n341 3.947
R614 VP.n747 VP.n746 3.588
R615 VP.n744 VP.n741 3.588
R616 VP.n678 VP.n677 3.588
R617 VP.n675 VP.n672 3.588
R618 VP.n609 VP.n608 3.588
R619 VP.n606 VP.n603 3.588
R620 VP.n539 VP.n538 3.588
R621 VP.n536 VP.n533 3.588
R622 VP.n470 VP.n469 3.588
R623 VP.n467 VP.n464 3.588
R624 VP.n119 VP.n118 3.588
R625 VP.n116 VP.n113 3.588
R626 VP.n50 VP.n49 3.588
R627 VP.n47 VP.n44 3.588
R628 VP.n258 VP.n257 3.588
R629 VP.n255 VP.n252 3.588
R630 VP.n189 VP.n188 3.588
R631 VP.n186 VP.n183 3.588
R632 VP.n397 VP.n396 3.588
R633 VP.n394 VP.n391 3.588
R634 VP.n328 VP.n327 3.588
R635 VP.n325 VP.n322 3.588
R636 VP.n708 VP.n707 3.396
R637 VP.n754 VP.n753 3.229
R638 VP.n753 VP.n752 3.229
R639 VP.n685 VP.n684 3.229
R640 VP.n684 VP.n683 3.229
R641 VP.n616 VP.n615 3.229
R642 VP.n615 VP.n614 3.229
R643 VP.n546 VP.n545 3.229
R644 VP.n545 VP.n544 3.229
R645 VP.n477 VP.n476 3.229
R646 VP.n476 VP.n475 3.229
R647 VP.n126 VP.n125 3.229
R648 VP.n125 VP.n124 3.229
R649 VP.n57 VP.n56 3.229
R650 VP.n56 VP.n55 3.229
R651 VP.n265 VP.n264 3.229
R652 VP.n264 VP.n263 3.229
R653 VP.n196 VP.n195 3.229
R654 VP.n195 VP.n194 3.229
R655 VP.n404 VP.n403 3.229
R656 VP.n403 VP.n402 3.229
R657 VP.n335 VP.n334 3.229
R658 VP.n334 VP.n333 3.229
R659 VP.n431 VP.n430 3.177
R660 VP.n289 VP.n288 3.177
R661 VP.n639 VP.n638 2.984
R662 VP.n570 VP.n569 2.984
R663 VP.n500 VP.n499 2.984
R664 VP.n80 VP.n79 2.984
R665 VP.n11 VP.n10 2.984
R666 VP.n219 VP.n218 2.984
R667 VP.n150 VP.n149 2.984
R668 VP.n358 VP.n357 2.984
R669 VP.n755 VP.n754 2.87
R670 VP.n752 VP.n749 2.87
R671 VP.n686 VP.n685 2.87
R672 VP.n683 VP.n680 2.87
R673 VP.n617 VP.n616 2.87
R674 VP.n614 VP.n611 2.87
R675 VP.n547 VP.n546 2.87
R676 VP.n544 VP.n541 2.87
R677 VP.n478 VP.n477 2.87
R678 VP.n475 VP.n472 2.87
R679 VP.n127 VP.n126 2.87
R680 VP.n124 VP.n121 2.87
R681 VP.n58 VP.n57 2.87
R682 VP.n55 VP.n52 2.87
R683 VP.n266 VP.n265 2.87
R684 VP.n263 VP.n260 2.87
R685 VP.n197 VP.n196 2.87
R686 VP.n194 VP.n191 2.87
R687 VP.n405 VP.n404 2.87
R688 VP.n402 VP.n399 2.87
R689 VP.n336 VP.n335 2.87
R690 VP.n333 VP.n330 2.87
R691 VP.n746 VP.n745 2.511
R692 VP.n745 VP.n744 2.511
R693 VP.n677 VP.n676 2.511
R694 VP.n676 VP.n675 2.511
R695 VP.n608 VP.n607 2.511
R696 VP.n607 VP.n606 2.511
R697 VP.n538 VP.n537 2.511
R698 VP.n537 VP.n536 2.511
R699 VP.n469 VP.n468 2.511
R700 VP.n468 VP.n467 2.511
R701 VP.n118 VP.n117 2.511
R702 VP.n117 VP.n116 2.511
R703 VP.n49 VP.n48 2.511
R704 VP.n48 VP.n47 2.511
R705 VP.n257 VP.n256 2.511
R706 VP.n256 VP.n255 2.511
R707 VP.n188 VP.n187 2.511
R708 VP.n187 VP.n186 2.511
R709 VP.n396 VP.n395 2.511
R710 VP.n395 VP.n394 2.511
R711 VP.n327 VP.n326 2.511
R712 VP.n326 VP.n325 2.511
R713 VP.n763 VP.n762 2.152
R714 VP.n760 VP.n757 2.152
R715 VP.n694 VP.n693 2.152
R716 VP.n691 VP.n688 2.152
R717 VP.n625 VP.n624 2.152
R718 VP.n622 VP.n619 2.152
R719 VP.n555 VP.n554 2.152
R720 VP.n552 VP.n549 2.152
R721 VP.n486 VP.n485 2.152
R722 VP.n483 VP.n480 2.152
R723 VP.n135 VP.n134 2.152
R724 VP.n132 VP.n129 2.152
R725 VP.n66 VP.n65 2.152
R726 VP.n63 VP.n60 2.152
R727 VP.n274 VP.n273 2.152
R728 VP.n271 VP.n268 2.152
R729 VP.n205 VP.n204 2.152
R730 VP.n202 VP.n199 2.152
R731 VP.n413 VP.n412 2.152
R732 VP.n410 VP.n407 2.152
R733 VP.n344 VP.n343 2.152
R734 VP.n341 VP.n338 2.152
R735 VP.n738 VP.n737 1.794
R736 VP.n737 VP.n736 1.794
R737 VP.n669 VP.n668 1.794
R738 VP.n668 VP.n667 1.794
R739 VP.n600 VP.n599 1.794
R740 VP.n599 VP.n598 1.794
R741 VP.n530 VP.n529 1.794
R742 VP.n529 VP.n528 1.794
R743 VP.n461 VP.n460 1.794
R744 VP.n460 VP.n459 1.794
R745 VP.n110 VP.n109 1.794
R746 VP.n109 VP.n108 1.794
R747 VP.n41 VP.n40 1.794
R748 VP.n40 VP.n39 1.794
R749 VP.n249 VP.n248 1.794
R750 VP.n248 VP.n247 1.794
R751 VP.n180 VP.n179 1.794
R752 VP.n179 VP.n178 1.794
R753 VP.n388 VP.n387 1.794
R754 VP.n387 VP.n386 1.794
R755 VP.n319 VP.n318 1.794
R756 VP.n318 VP.n317 1.794
R757 VP.n698 VP.n697 1.076
R758 VP.n701 VP.n698 1.076
R759 VP.n629 VP.n628 1.076
R760 VP.n632 VP.n629 1.076
R761 VP.n560 VP.n559 1.076
R762 VP.n563 VP.n560 1.076
R763 VP.n490 VP.n489 1.076
R764 VP.n493 VP.n490 1.076
R765 VP.n421 VP.n420 1.076
R766 VP.n424 VP.n421 1.076
R767 VP.n70 VP.n69 1.076
R768 VP.n73 VP.n70 1.076
R769 VP.n1 VP.n0 1.076
R770 VP.n4 VP.n1 1.076
R771 VP.n209 VP.n208 1.076
R772 VP.n212 VP.n209 1.076
R773 VP.n140 VP.n139 1.076
R774 VP.n143 VP.n140 1.076
R775 VP.n348 VP.n347 1.076
R776 VP.n351 VP.n348 1.076
R777 VP.n279 VP.n278 1.076
R778 VP.n282 VP.n279 1.076
R779 VP.n418 VP.n417 0.491
R780 VP.n419 VP.n418 0.483
R781 VP.n706 VP.n705 0.358
R782 VP.n709 VP.n706 0.358
R783 VP.n637 VP.n636 0.358
R784 VP.n640 VP.n637 0.358
R785 VP.n568 VP.n567 0.358
R786 VP.n571 VP.n568 0.358
R787 VP.n498 VP.n497 0.358
R788 VP.n501 VP.n498 0.358
R789 VP.n429 VP.n428 0.358
R790 VP.n432 VP.n429 0.358
R791 VP.n78 VP.n77 0.358
R792 VP.n81 VP.n78 0.358
R793 VP.n9 VP.n8 0.358
R794 VP.n12 VP.n9 0.358
R795 VP.n217 VP.n216 0.358
R796 VP.n220 VP.n217 0.358
R797 VP.n148 VP.n147 0.358
R798 VP.n151 VP.n148 0.358
R799 VP.n356 VP.n355 0.358
R800 VP.n359 VP.n356 0.358
R801 VP.n287 VP.n286 0.358
R802 VP.n290 VP.n287 0.358
R803 VP VP.n769 0.341
R804 VP.n728 VP.n727 0.144
R805 VP.n725 VP.n724 0.144
R806 VP.n722 VP.n721 0.144
R807 VP.n719 VP.n718 0.144
R808 VP.n716 VP.n715 0.144
R809 VP.n659 VP.n658 0.144
R810 VP.n656 VP.n655 0.144
R811 VP.n653 VP.n652 0.144
R812 VP.n650 VP.n649 0.144
R813 VP.n647 VP.n646 0.144
R814 VP.n590 VP.n589 0.144
R815 VP.n587 VP.n586 0.144
R816 VP.n584 VP.n583 0.144
R817 VP.n581 VP.n580 0.144
R818 VP.n578 VP.n577 0.144
R819 VP.n520 VP.n519 0.144
R820 VP.n517 VP.n516 0.144
R821 VP.n514 VP.n513 0.144
R822 VP.n511 VP.n510 0.144
R823 VP.n508 VP.n507 0.144
R824 VP.n451 VP.n450 0.144
R825 VP.n448 VP.n447 0.144
R826 VP.n445 VP.n444 0.144
R827 VP.n442 VP.n441 0.144
R828 VP.n439 VP.n438 0.144
R829 VP.n100 VP.n99 0.144
R830 VP.n97 VP.n96 0.144
R831 VP.n94 VP.n93 0.144
R832 VP.n91 VP.n90 0.144
R833 VP.n88 VP.n87 0.144
R834 VP.n31 VP.n30 0.144
R835 VP.n28 VP.n27 0.144
R836 VP.n25 VP.n24 0.144
R837 VP.n22 VP.n21 0.144
R838 VP.n19 VP.n18 0.144
R839 VP.n239 VP.n238 0.144
R840 VP.n236 VP.n235 0.144
R841 VP.n233 VP.n232 0.144
R842 VP.n230 VP.n229 0.144
R843 VP.n227 VP.n226 0.144
R844 VP.n170 VP.n169 0.144
R845 VP.n167 VP.n166 0.144
R846 VP.n164 VP.n163 0.144
R847 VP.n161 VP.n160 0.144
R848 VP.n158 VP.n157 0.144
R849 VP.n378 VP.n377 0.144
R850 VP.n375 VP.n374 0.144
R851 VP.n372 VP.n371 0.144
R852 VP.n369 VP.n368 0.144
R853 VP.n366 VP.n365 0.144
R854 VP.n309 VP.n308 0.144
R855 VP.n306 VP.n305 0.144
R856 VP.n303 VP.n302 0.144
R857 VP.n300 VP.n299 0.144
R858 VP.n297 VP.n296 0.144
R859 VP VP.n419 0.124
R860 VP.n715 VP.n714 0.043
R861 VP.n646 VP.n645 0.043
R862 VP.n577 VP.n576 0.043
R863 VP.n507 VP.n506 0.043
R864 VP.n438 VP.n437 0.043
R865 VP.n87 VP.n86 0.043
R866 VP.n18 VP.n17 0.043
R867 VP.n226 VP.n225 0.043
R868 VP.n157 VP.n156 0.043
R869 VP.n365 VP.n364 0.043
R870 VP.n296 VP.n295 0.043
R871 VP.n718 VP.n717 0.038
R872 VP.n649 VP.n648 0.038
R873 VP.n580 VP.n579 0.038
R874 VP.n510 VP.n509 0.038
R875 VP.n441 VP.n440 0.038
R876 VP.n90 VP.n89 0.038
R877 VP.n21 VP.n20 0.038
R878 VP.n229 VP.n228 0.038
R879 VP.n160 VP.n159 0.038
R880 VP.n368 VP.n367 0.038
R881 VP.n299 VP.n298 0.038
R882 VP.n721 VP.n720 0.032
R883 VP.n652 VP.n651 0.032
R884 VP.n583 VP.n582 0.032
R885 VP.n513 VP.n512 0.032
R886 VP.n444 VP.n443 0.032
R887 VP.n93 VP.n92 0.032
R888 VP.n24 VP.n23 0.032
R889 VP.n232 VP.n231 0.032
R890 VP.n163 VP.n162 0.032
R891 VP.n371 VP.n370 0.032
R892 VP.n302 VP.n301 0.032
R893 VP.n729 VP.n728 0.029
R894 VP.n660 VP.n659 0.029
R895 VP.n591 VP.n590 0.029
R896 VP.n521 VP.n520 0.029
R897 VP.n452 VP.n451 0.029
R898 VP.n101 VP.n100 0.029
R899 VP.n32 VP.n31 0.029
R900 VP.n240 VP.n239 0.029
R901 VP.n171 VP.n170 0.029
R902 VP.n379 VP.n378 0.029
R903 VP.n310 VP.n309 0.029
R904 VP.n724 VP.n723 0.027
R905 VP.n655 VP.n654 0.027
R906 VP.n586 VP.n585 0.027
R907 VP.n516 VP.n515 0.027
R908 VP.n447 VP.n446 0.027
R909 VP.n96 VP.n95 0.027
R910 VP.n27 VP.n26 0.027
R911 VP.n235 VP.n234 0.027
R912 VP.n166 VP.n165 0.027
R913 VP.n374 VP.n373 0.027
R914 VP.n305 VP.n304 0.027
R915 VP.n726 VP.n725 0.024
R916 VP.n657 VP.n656 0.024
R917 VP.n588 VP.n587 0.024
R918 VP.n518 VP.n517 0.024
R919 VP.n449 VP.n448 0.024
R920 VP.n98 VP.n97 0.024
R921 VP.n29 VP.n28 0.024
R922 VP.n237 VP.n236 0.024
R923 VP.n168 VP.n167 0.024
R924 VP.n376 VP.n375 0.024
R925 VP.n307 VP.n306 0.024
R926 VP.n727 VP.n726 0.021
R927 VP.n658 VP.n657 0.021
R928 VP.n589 VP.n588 0.021
R929 VP.n519 VP.n518 0.021
R930 VP.n450 VP.n449 0.021
R931 VP.n99 VP.n98 0.021
R932 VP.n30 VP.n29 0.021
R933 VP.n238 VP.n237 0.021
R934 VP.n169 VP.n168 0.021
R935 VP.n377 VP.n376 0.021
R936 VP.n308 VP.n307 0.021
R937 VP.n723 VP.n722 0.019
R938 VP.n654 VP.n653 0.019
R939 VP.n585 VP.n584 0.019
R940 VP.n515 VP.n514 0.019
R941 VP.n446 VP.n445 0.019
R942 VP.n95 VP.n94 0.019
R943 VP.n26 VP.n25 0.019
R944 VP.n234 VP.n233 0.019
R945 VP.n165 VP.n164 0.019
R946 VP.n373 VP.n372 0.019
R947 VP.n304 VP.n303 0.019
R948 VP.n730 VP.n729 0.016
R949 VP.n661 VP.n660 0.016
R950 VP.n592 VP.n591 0.016
R951 VP.n522 VP.n521 0.016
R952 VP.n453 VP.n452 0.016
R953 VP.n102 VP.n101 0.016
R954 VP.n33 VP.n32 0.016
R955 VP.n241 VP.n240 0.016
R956 VP.n172 VP.n171 0.016
R957 VP.n380 VP.n379 0.016
R958 VP.n311 VP.n310 0.016
R959 VP.n720 VP.n719 0.013
R960 VP.n651 VP.n650 0.013
R961 VP.n582 VP.n581 0.013
R962 VP.n512 VP.n511 0.013
R963 VP.n443 VP.n442 0.013
R964 VP.n92 VP.n91 0.013
R965 VP.n23 VP.n22 0.013
R966 VP.n231 VP.n230 0.013
R967 VP.n162 VP.n161 0.013
R968 VP.n370 VP.n369 0.013
R969 VP.n301 VP.n300 0.013
R970 VP.n717 VP.n716 0.008
R971 VP.n648 VP.n647 0.008
R972 VP.n579 VP.n578 0.008
R973 VP.n509 VP.n508 0.008
R974 VP.n440 VP.n439 0.008
R975 VP.n89 VP.n88 0.008
R976 VP.n20 VP.n19 0.008
R977 VP.n228 VP.n227 0.008
R978 VP.n159 VP.n158 0.008
R979 VP.n367 VP.n366 0.008
R980 VP.n298 VP.n297 0.008
R981 VP.n714 VP.n713 0.002
R982 VP.n645 VP.n644 0.002
R983 VP.n576 VP.n575 0.002
R984 VP.n506 VP.n505 0.002
R985 VP.n437 VP.n436 0.002
R986 VP.n86 VP.n85 0.002
R987 VP.n17 VP.n16 0.002
R988 VP.n225 VP.n224 0.002
R989 VP.n156 VP.n155 0.002
R990 VP.n364 VP.n363 0.002
R991 VP.n295 VP.n294 0.002
R992 a_6260_5590.n144 a_6260_5590.n143 287.957
R993 a_6260_5590.n143 a_6260_5590.n142 186.836
R994 a_6260_5590.n143 a_6260_5590.n75 169.426
R995 a_6260_5590.n91 a_6260_5590.t0 64.755
R996 a_6260_5590.n24 a_6260_5590.t1 64.755
R997 a_6260_5590.t2 a_6260_5590.n199 53.727
R998 a_6260_5590.n142 a_6260_5590.n107 49.503
R999 a_6260_5590.n75 a_6260_5590.n40 49.503
R1000 a_6260_5590.n145 a_6260_5590.n144 49.503
R1001 a_6260_5590.n136 a_6260_5590.n135 32.833
R1002 a_6260_5590.n69 a_6260_5590.n68 32.833
R1003 a_6260_5590.n3 a_6260_5590.n2 32.833
R1004 a_6260_5590.n25 a_6260_5590.n24 30.598
R1005 a_6260_5590.n92 a_6260_5590.n91 30.598
R1006 a_6260_5590.t2 a_6260_5590.n159 95.496
R1007 a_6260_5590.n128 a_6260_5590.n127 26.863
R1008 a_6260_5590.n61 a_6260_5590.n60 26.863
R1009 a_6260_5590.n164 a_6260_5590.n163 26.863
R1010 a_6260_5590.n120 a_6260_5590.n119 20.893
R1011 a_6260_5590.n53 a_6260_5590.n52 20.893
R1012 a_6260_5590.n172 a_6260_5590.n171 20.893
R1013 a_6260_5590.n88 a_6260_5590.n87 15
R1014 a_6260_5590.n80 a_6260_5590.n79 15
R1015 a_6260_5590.n113 a_6260_5590.n112 15
R1016 a_6260_5590.n121 a_6260_5590.n120 15
R1017 a_6260_5590.n129 a_6260_5590.n128 15
R1018 a_6260_5590.n90 a_6260_5590.n89 15
R1019 a_6260_5590.n82 a_6260_5590.n81 15
R1020 a_6260_5590.n110 a_6260_5590.n109 15
R1021 a_6260_5590.n118 a_6260_5590.n117 15
R1022 a_6260_5590.n126 a_6260_5590.n125 15
R1023 a_6260_5590.n134 a_6260_5590.n133 15
R1024 a_6260_5590.n137 a_6260_5590.n136 15
R1025 a_6260_5590.n21 a_6260_5590.n20 15
R1026 a_6260_5590.n13 a_6260_5590.n12 15
R1027 a_6260_5590.n46 a_6260_5590.n45 15
R1028 a_6260_5590.n54 a_6260_5590.n53 15
R1029 a_6260_5590.n62 a_6260_5590.n61 15
R1030 a_6260_5590.n70 a_6260_5590.n69 15
R1031 a_6260_5590.n23 a_6260_5590.n22 15
R1032 a_6260_5590.n15 a_6260_5590.n14 15
R1033 a_6260_5590.n43 a_6260_5590.n42 15
R1034 a_6260_5590.n51 a_6260_5590.n50 15
R1035 a_6260_5590.n59 a_6260_5590.n58 15
R1036 a_6260_5590.n67 a_6260_5590.n66 15
R1037 a_6260_5590.n197 a_6260_5590.n196 15
R1038 a_6260_5590.n189 a_6260_5590.n188 15
R1039 a_6260_5590.n181 a_6260_5590.n180 15
R1040 a_6260_5590.n173 a_6260_5590.n172 15
R1041 a_6260_5590.n165 a_6260_5590.n164 15
R1042 a_6260_5590.n199 a_6260_5590.n198 15
R1043 a_6260_5590.n191 a_6260_5590.n190 15
R1044 a_6260_5590.n183 a_6260_5590.n182 15
R1045 a_6260_5590.n175 a_6260_5590.n174 15
R1046 a_6260_5590.n167 a_6260_5590.n166 15
R1047 a_6260_5590.n1 a_6260_5590.n0 15
R1048 a_6260_5590.n4 a_6260_5590.n3 15
R1049 a_6260_5590.n112 a_6260_5590.n111 14.924
R1050 a_6260_5590.n45 a_6260_5590.n44 14.924
R1051 a_6260_5590.n180 a_6260_5590.n179 14.924
R1052 a_6260_5590.n91 a_6260_5590.n90 14.123
R1053 a_6260_5590.n24 a_6260_5590.n23 14.123
R1054 a_6260_5590.n141 a_6260_5590.n140 13.544
R1055 a_6260_5590.n74 a_6260_5590.n73 13.544
R1056 a_6260_5590.n8 a_6260_5590.n7 13.544
R1057 a_6260_5590.n83 a_6260_5590.n82 12.917
R1058 a_6260_5590.n110 a_6260_5590.n108 12.917
R1059 a_6260_5590.n118 a_6260_5590.n116 12.917
R1060 a_6260_5590.n126 a_6260_5590.n124 12.917
R1061 a_6260_5590.n134 a_6260_5590.n132 12.917
R1062 a_6260_5590.n67 a_6260_5590.n65 12.917
R1063 a_6260_5590.n59 a_6260_5590.n57 12.917
R1064 a_6260_5590.n51 a_6260_5590.n49 12.917
R1065 a_6260_5590.n43 a_6260_5590.n41 12.917
R1066 a_6260_5590.n16 a_6260_5590.n15 12.917
R1067 a_6260_5590.n192 a_6260_5590.n191 12.917
R1068 a_6260_5590.n184 a_6260_5590.n183 12.917
R1069 a_6260_5590.n176 a_6260_5590.n175 12.917
R1070 a_6260_5590.n168 a_6260_5590.n167 12.917
R1071 a_6260_5590.n79 a_6260_5590.n78 8.954
R1072 a_6260_5590.n12 a_6260_5590.n11 8.954
R1073 a_6260_5590.n188 a_6260_5590.n187 8.954
R1074 a_6260_5590.n142 a_6260_5590.n141 8.805
R1075 a_6260_5590.n75 a_6260_5590.n74 8.805
R1076 a_6260_5590.n144 a_6260_5590.n8 8.805
R1077 a_6260_5590.n90 a_6260_5590.n88 5.741
R1078 a_6260_5590.n84 a_6260_5590.n83 5.741
R1079 a_6260_5590.n17 a_6260_5590.n16 5.741
R1080 a_6260_5590.n23 a_6260_5590.n21 5.741
R1081 a_6260_5590.n198 a_6260_5590.n197 5.741
R1082 a_6260_5590.n193 a_6260_5590.n192 5.741
R1083 a_6260_5590.n82 a_6260_5590.n80 5.023
R1084 a_6260_5590.n15 a_6260_5590.n13 5.023
R1085 a_6260_5590.n191 a_6260_5590.n189 5.023
R1086 a_6260_5590.n185 a_6260_5590.n184 5.023
R1087 a_6260_5590.n113 a_6260_5590.n110 4.305
R1088 a_6260_5590.n116 a_6260_5590.n115 4.305
R1089 a_6260_5590.n49 a_6260_5590.n48 4.305
R1090 a_6260_5590.n46 a_6260_5590.n43 4.305
R1091 a_6260_5590.n183 a_6260_5590.n181 4.305
R1092 a_6260_5590.n177 a_6260_5590.n176 4.305
R1093 a_6260_5590.n138 a_6260_5590.n137 3.947
R1094 a_6260_5590.n139 a_6260_5590.n138 3.947
R1095 a_6260_5590.n72 a_6260_5590.n71 3.947
R1096 a_6260_5590.n71 a_6260_5590.n70 3.947
R1097 a_6260_5590.n5 a_6260_5590.n4 3.947
R1098 a_6260_5590.n6 a_6260_5590.n5 3.947
R1099 a_6260_5590.n121 a_6260_5590.n118 3.588
R1100 a_6260_5590.n124 a_6260_5590.n123 3.588
R1101 a_6260_5590.n57 a_6260_5590.n56 3.588
R1102 a_6260_5590.n54 a_6260_5590.n51 3.588
R1103 a_6260_5590.n175 a_6260_5590.n173 3.588
R1104 a_6260_5590.n169 a_6260_5590.n168 3.588
R1105 a_6260_5590.n130 a_6260_5590.n129 3.229
R1106 a_6260_5590.n131 a_6260_5590.n130 3.229
R1107 a_6260_5590.n64 a_6260_5590.n63 3.229
R1108 a_6260_5590.n63 a_6260_5590.n62 3.229
R1109 a_6260_5590.n165 a_6260_5590.n162 3.229
R1110 a_6260_5590.n162 a_6260_5590.n161 3.229
R1111 a_6260_5590.n87 a_6260_5590.n86 2.984
R1112 a_6260_5590.n20 a_6260_5590.n19 2.984
R1113 a_6260_5590.n196 a_6260_5590.n195 2.984
R1114 a_6260_5590.n129 a_6260_5590.n126 2.87
R1115 a_6260_5590.n132 a_6260_5590.n131 2.87
R1116 a_6260_5590.n65 a_6260_5590.n64 2.87
R1117 a_6260_5590.n62 a_6260_5590.n59 2.87
R1118 a_6260_5590.n167 a_6260_5590.n165 2.87
R1119 a_6260_5590.n161 a_6260_5590.n160 2.87
R1120 a_6260_5590.n122 a_6260_5590.n121 2.511
R1121 a_6260_5590.n123 a_6260_5590.n122 2.511
R1122 a_6260_5590.n56 a_6260_5590.n55 2.511
R1123 a_6260_5590.n55 a_6260_5590.n54 2.511
R1124 a_6260_5590.n173 a_6260_5590.n170 2.511
R1125 a_6260_5590.n170 a_6260_5590.n169 2.511
R1126 a_6260_5590.n137 a_6260_5590.n134 2.152
R1127 a_6260_5590.n140 a_6260_5590.n139 2.152
R1128 a_6260_5590.n73 a_6260_5590.n72 2.152
R1129 a_6260_5590.n70 a_6260_5590.n67 2.152
R1130 a_6260_5590.n4 a_6260_5590.n1 2.152
R1131 a_6260_5590.n7 a_6260_5590.n6 2.152
R1132 a_6260_5590.n114 a_6260_5590.n113 1.794
R1133 a_6260_5590.n115 a_6260_5590.n114 1.794
R1134 a_6260_5590.n48 a_6260_5590.n47 1.794
R1135 a_6260_5590.n47 a_6260_5590.n46 1.794
R1136 a_6260_5590.n181 a_6260_5590.n178 1.794
R1137 a_6260_5590.n178 a_6260_5590.n177 1.794
R1138 a_6260_5590.n80 a_6260_5590.n77 1.076
R1139 a_6260_5590.n77 a_6260_5590.n76 1.076
R1140 a_6260_5590.n10 a_6260_5590.n9 1.076
R1141 a_6260_5590.n13 a_6260_5590.n10 1.076
R1142 a_6260_5590.n189 a_6260_5590.n186 1.076
R1143 a_6260_5590.n186 a_6260_5590.n185 1.076
R1144 a_6260_5590.n88 a_6260_5590.n85 0.358
R1145 a_6260_5590.n85 a_6260_5590.n84 0.358
R1146 a_6260_5590.n18 a_6260_5590.n17 0.358
R1147 a_6260_5590.n21 a_6260_5590.n18 0.358
R1148 a_6260_5590.n197 a_6260_5590.n194 0.358
R1149 a_6260_5590.n194 a_6260_5590.n193 0.358
R1150 a_6260_5590.n93 a_6260_5590.n92 0.144
R1151 a_6260_5590.n96 a_6260_5590.n95 0.144
R1152 a_6260_5590.n99 a_6260_5590.n98 0.144
R1153 a_6260_5590.n102 a_6260_5590.n101 0.144
R1154 a_6260_5590.n105 a_6260_5590.n104 0.144
R1155 a_6260_5590.n38 a_6260_5590.n37 0.144
R1156 a_6260_5590.n35 a_6260_5590.n34 0.144
R1157 a_6260_5590.n32 a_6260_5590.n31 0.144
R1158 a_6260_5590.n29 a_6260_5590.n28 0.144
R1159 a_6260_5590.n26 a_6260_5590.n25 0.144
R1160 a_6260_5590.n157 a_6260_5590.n156 0.144
R1161 a_6260_5590.n154 a_6260_5590.n153 0.144
R1162 a_6260_5590.n151 a_6260_5590.n150 0.144
R1163 a_6260_5590.n148 a_6260_5590.n147 0.144
R1164 a_6260_5590.n95 a_6260_5590.n94 0.038
R1165 a_6260_5590.n28 a_6260_5590.n27 0.038
R1166 a_6260_5590.n158 a_6260_5590.n157 0.038
R1167 a_6260_5590.n98 a_6260_5590.n97 0.032
R1168 a_6260_5590.n31 a_6260_5590.n30 0.032
R1169 a_6260_5590.n155 a_6260_5590.n154 0.032
R1170 a_6260_5590.n106 a_6260_5590.n105 0.029
R1171 a_6260_5590.n39 a_6260_5590.n38 0.029
R1172 a_6260_5590.n147 a_6260_5590.n146 0.029
R1173 a_6260_5590.n101 a_6260_5590.n100 0.027
R1174 a_6260_5590.n34 a_6260_5590.n33 0.027
R1175 a_6260_5590.n152 a_6260_5590.n151 0.027
R1176 a_6260_5590.n103 a_6260_5590.n102 0.024
R1177 a_6260_5590.n36 a_6260_5590.n35 0.024
R1178 a_6260_5590.n150 a_6260_5590.n149 0.024
R1179 a_6260_5590.n104 a_6260_5590.n103 0.021
R1180 a_6260_5590.n37 a_6260_5590.n36 0.021
R1181 a_6260_5590.n149 a_6260_5590.n148 0.021
R1182 a_6260_5590.n100 a_6260_5590.n99 0.019
R1183 a_6260_5590.n33 a_6260_5590.n32 0.019
R1184 a_6260_5590.n153 a_6260_5590.n152 0.019
R1185 a_6260_5590.n107 a_6260_5590.n106 0.016
R1186 a_6260_5590.n40 a_6260_5590.n39 0.016
R1187 a_6260_5590.n146 a_6260_5590.n145 0.016
R1188 a_6260_5590.n97 a_6260_5590.n96 0.013
R1189 a_6260_5590.n30 a_6260_5590.n29 0.013
R1190 a_6260_5590.n156 a_6260_5590.n155 0.013
R1191 a_6260_5590.n94 a_6260_5590.n93 0.008
R1192 a_6260_5590.n27 a_6260_5590.n26 0.008
R1193 a_6260_5590.n159 a_6260_5590.n158 0.008
R1194 VCT.n74 VCT.t5 1306.2
R1195 VCT.n63 VCT.n62 1060.4
R1196 VCT.n49 VCT.t1 1060.4
R1197 VCT.n35 VCT.n34 1060.4
R1198 VCT.n21 VCT.n20 1060.4
R1199 VCT.n7 VCT.n6 1060.4
R1200 VCT.n63 VCT.n61 906.159
R1201 VCT.n64 VCT.n60 906.159
R1202 VCT.n65 VCT.n59 906.159
R1203 VCT.n66 VCT.t4 906.159
R1204 VCT.n67 VCT.n58 906.159
R1205 VCT.n68 VCT.n57 906.159
R1206 VCT.n69 VCT.n56 906.159
R1207 VCT.n49 VCT.n48 906.159
R1208 VCT.n50 VCT.n47 906.159
R1209 VCT.n51 VCT.n46 906.159
R1210 VCT.n52 VCT.n45 906.159
R1211 VCT.n53 VCT.n44 906.159
R1212 VCT.n54 VCT.n43 906.159
R1213 VCT.n55 VCT.n42 906.159
R1214 VCT.n35 VCT.n33 906.159
R1215 VCT.n36 VCT.n32 906.159
R1216 VCT.n37 VCT.n31 906.159
R1217 VCT.n38 VCT.t3 906.159
R1218 VCT.n39 VCT.n30 906.159
R1219 VCT.n40 VCT.n29 906.159
R1220 VCT.n41 VCT.n28 906.159
R1221 VCT.n21 VCT.n19 906.159
R1222 VCT.n22 VCT.n18 906.159
R1223 VCT.n23 VCT.n17 906.159
R1224 VCT.n24 VCT.n16 906.159
R1225 VCT.n25 VCT.t0 906.159
R1226 VCT.n26 VCT.n15 906.159
R1227 VCT.n27 VCT.n14 906.159
R1228 VCT.n7 VCT.n5 906.159
R1229 VCT.n8 VCT.n4 906.159
R1230 VCT.n9 VCT.n3 906.159
R1231 VCT.n10 VCT.n2 906.159
R1232 VCT.n11 VCT.n1 906.159
R1233 VCT.n12 VCT.n0 906.159
R1234 VCT.n13 VCT.t2 906.159
R1235 VCT.n70 VCT.n69 252.567
R1236 VCT.n72 VCT.n27 251.031
R1237 VCT.n70 VCT.n55 251.027
R1238 VCT.n71 VCT.n41 250.916
R1239 VCT.n73 VCT.n13 250.756
R1240 VCT.n68 VCT.n67 154.24
R1241 VCT.n67 VCT.n66 154.24
R1242 VCT.n66 VCT.n65 154.24
R1243 VCT.n65 VCT.n64 154.24
R1244 VCT.n64 VCT.n63 154.24
R1245 VCT.n54 VCT.n53 154.24
R1246 VCT.n53 VCT.n52 154.24
R1247 VCT.n52 VCT.n51 154.24
R1248 VCT.n51 VCT.n50 154.24
R1249 VCT.n50 VCT.n49 154.24
R1250 VCT.n40 VCT.n39 154.24
R1251 VCT.n39 VCT.n38 154.24
R1252 VCT.n38 VCT.n37 154.24
R1253 VCT.n37 VCT.n36 154.24
R1254 VCT.n36 VCT.n35 154.24
R1255 VCT.n26 VCT.n25 154.24
R1256 VCT.n25 VCT.n24 154.24
R1257 VCT.n24 VCT.n23 154.24
R1258 VCT.n23 VCT.n22 154.24
R1259 VCT.n22 VCT.n21 154.24
R1260 VCT.n12 VCT.n11 154.24
R1261 VCT.n11 VCT.n10 154.24
R1262 VCT.n10 VCT.n9 154.24
R1263 VCT.n9 VCT.n8 154.24
R1264 VCT.n8 VCT.n7 154.24
R1265 VCT.n69 VCT.n68 148.215
R1266 VCT.n55 VCT.n54 148.215
R1267 VCT.n41 VCT.n40 148.215
R1268 VCT.n27 VCT.n26 148.215
R1269 VCT.n13 VCT.n12 148.215
R1270 VCT.n74 VCT.n73 3.776
R1271 VCT VCT.n74 2.199
R1272 VCT.n72 VCT.n71 1.789
R1273 VCT.n71 VCT.n70 1.694
R1274 VCT.n73 VCT.n72 1.59
R1275 a_9348_5588.n143 a_9348_5588.n75 238.293
R1276 a_9348_5588.n143 a_9348_5588.n142 186.678
R1277 a_9348_5588.n144 a_9348_5588.n143 160.08
R1278 a_9348_5588.n24 a_9348_5588.t2 68.375
R1279 a_9348_5588.n91 a_9348_5588.t1 64.755
R1280 a_9348_5588.t0 a_9348_5588.n199 53.727
R1281 a_9348_5588.n142 a_9348_5588.n107 49.503
R1282 a_9348_5588.n75 a_9348_5588.n40 49.503
R1283 a_9348_5588.n145 a_9348_5588.n144 49.503
R1284 a_9348_5588.n69 a_9348_5588.n68 34.951
R1285 a_9348_5588.n136 a_9348_5588.n135 32.833
R1286 a_9348_5588.n3 a_9348_5588.n2 32.833
R1287 a_9348_5588.n25 a_9348_5588.n24 30.732
R1288 a_9348_5588.n92 a_9348_5588.n91 30.598
R1289 a_9348_5588.t0 a_9348_5588.n159 95.496
R1290 a_9348_5588.n61 a_9348_5588.n60 28.596
R1291 a_9348_5588.n128 a_9348_5588.n127 26.863
R1292 a_9348_5588.n164 a_9348_5588.n163 26.863
R1293 a_9348_5588.n53 a_9348_5588.n52 22.241
R1294 a_9348_5588.n120 a_9348_5588.n119 20.893
R1295 a_9348_5588.n172 a_9348_5588.n171 20.893
R1296 a_9348_5588.n45 a_9348_5588.n44 15.887
R1297 a_9348_5588.n88 a_9348_5588.n87 15
R1298 a_9348_5588.n80 a_9348_5588.n79 15
R1299 a_9348_5588.n113 a_9348_5588.n112 15
R1300 a_9348_5588.n121 a_9348_5588.n120 15
R1301 a_9348_5588.n129 a_9348_5588.n128 15
R1302 a_9348_5588.n90 a_9348_5588.n89 15
R1303 a_9348_5588.n82 a_9348_5588.n81 15
R1304 a_9348_5588.n110 a_9348_5588.n109 15
R1305 a_9348_5588.n118 a_9348_5588.n117 15
R1306 a_9348_5588.n126 a_9348_5588.n125 15
R1307 a_9348_5588.n134 a_9348_5588.n133 15
R1308 a_9348_5588.n137 a_9348_5588.n136 15
R1309 a_9348_5588.n21 a_9348_5588.n20 15
R1310 a_9348_5588.n13 a_9348_5588.n12 15
R1311 a_9348_5588.n46 a_9348_5588.n45 15
R1312 a_9348_5588.n54 a_9348_5588.n53 15
R1313 a_9348_5588.n62 a_9348_5588.n61 15
R1314 a_9348_5588.n70 a_9348_5588.n69 15
R1315 a_9348_5588.n23 a_9348_5588.n22 15
R1316 a_9348_5588.n15 a_9348_5588.n14 15
R1317 a_9348_5588.n43 a_9348_5588.n42 15
R1318 a_9348_5588.n51 a_9348_5588.n50 15
R1319 a_9348_5588.n59 a_9348_5588.n58 15
R1320 a_9348_5588.n67 a_9348_5588.n66 15
R1321 a_9348_5588.n197 a_9348_5588.n196 15
R1322 a_9348_5588.n189 a_9348_5588.n188 15
R1323 a_9348_5588.n181 a_9348_5588.n180 15
R1324 a_9348_5588.n173 a_9348_5588.n172 15
R1325 a_9348_5588.n165 a_9348_5588.n164 15
R1326 a_9348_5588.n199 a_9348_5588.n198 15
R1327 a_9348_5588.n191 a_9348_5588.n190 15
R1328 a_9348_5588.n183 a_9348_5588.n182 15
R1329 a_9348_5588.n175 a_9348_5588.n174 15
R1330 a_9348_5588.n167 a_9348_5588.n166 15
R1331 a_9348_5588.n1 a_9348_5588.n0 15
R1332 a_9348_5588.n4 a_9348_5588.n3 15
R1333 a_9348_5588.n112 a_9348_5588.n111 14.924
R1334 a_9348_5588.n180 a_9348_5588.n179 14.924
R1335 a_9348_5588.n91 a_9348_5588.n90 14.123
R1336 a_9348_5588.n24 a_9348_5588.n23 14.071
R1337 a_9348_5588.n141 a_9348_5588.n140 13.544
R1338 a_9348_5588.n8 a_9348_5588.n7 13.544
R1339 a_9348_5588.n74 a_9348_5588.n73 13.532
R1340 a_9348_5588.n83 a_9348_5588.n82 12.917
R1341 a_9348_5588.n110 a_9348_5588.n108 12.917
R1342 a_9348_5588.n118 a_9348_5588.n116 12.917
R1343 a_9348_5588.n126 a_9348_5588.n124 12.917
R1344 a_9348_5588.n134 a_9348_5588.n132 12.917
R1345 a_9348_5588.n67 a_9348_5588.n65 12.917
R1346 a_9348_5588.n59 a_9348_5588.n57 12.917
R1347 a_9348_5588.n51 a_9348_5588.n49 12.917
R1348 a_9348_5588.n43 a_9348_5588.n41 12.917
R1349 a_9348_5588.n16 a_9348_5588.n15 12.917
R1350 a_9348_5588.n192 a_9348_5588.n191 12.917
R1351 a_9348_5588.n184 a_9348_5588.n183 12.917
R1352 a_9348_5588.n176 a_9348_5588.n175 12.917
R1353 a_9348_5588.n168 a_9348_5588.n167 12.917
R1354 a_9348_5588.n12 a_9348_5588.n11 9.532
R1355 a_9348_5588.n79 a_9348_5588.n78 8.954
R1356 a_9348_5588.n188 a_9348_5588.n187 8.954
R1357 a_9348_5588.n75 a_9348_5588.n74 8.82
R1358 a_9348_5588.n142 a_9348_5588.n141 8.805
R1359 a_9348_5588.n144 a_9348_5588.n8 8.805
R1360 a_9348_5588.n90 a_9348_5588.n88 5.741
R1361 a_9348_5588.n84 a_9348_5588.n83 5.741
R1362 a_9348_5588.n17 a_9348_5588.n16 5.741
R1363 a_9348_5588.n23 a_9348_5588.n21 5.741
R1364 a_9348_5588.n198 a_9348_5588.n197 5.741
R1365 a_9348_5588.n193 a_9348_5588.n192 5.741
R1366 a_9348_5588.n82 a_9348_5588.n80 5.023
R1367 a_9348_5588.n15 a_9348_5588.n13 5.023
R1368 a_9348_5588.n191 a_9348_5588.n189 5.023
R1369 a_9348_5588.n185 a_9348_5588.n184 5.023
R1370 a_9348_5588.n113 a_9348_5588.n110 4.305
R1371 a_9348_5588.n116 a_9348_5588.n115 4.305
R1372 a_9348_5588.n49 a_9348_5588.n48 4.305
R1373 a_9348_5588.n46 a_9348_5588.n43 4.305
R1374 a_9348_5588.n183 a_9348_5588.n181 4.305
R1375 a_9348_5588.n177 a_9348_5588.n176 4.305
R1376 a_9348_5588.n138 a_9348_5588.n137 3.947
R1377 a_9348_5588.n139 a_9348_5588.n138 3.947
R1378 a_9348_5588.n72 a_9348_5588.n71 3.947
R1379 a_9348_5588.n71 a_9348_5588.n70 3.947
R1380 a_9348_5588.n5 a_9348_5588.n4 3.947
R1381 a_9348_5588.n6 a_9348_5588.n5 3.947
R1382 a_9348_5588.n121 a_9348_5588.n118 3.588
R1383 a_9348_5588.n124 a_9348_5588.n123 3.588
R1384 a_9348_5588.n57 a_9348_5588.n56 3.588
R1385 a_9348_5588.n54 a_9348_5588.n51 3.588
R1386 a_9348_5588.n175 a_9348_5588.n173 3.588
R1387 a_9348_5588.n169 a_9348_5588.n168 3.588
R1388 a_9348_5588.n130 a_9348_5588.n129 3.229
R1389 a_9348_5588.n131 a_9348_5588.n130 3.229
R1390 a_9348_5588.n64 a_9348_5588.n63 3.229
R1391 a_9348_5588.n63 a_9348_5588.n62 3.229
R1392 a_9348_5588.n165 a_9348_5588.n162 3.229
R1393 a_9348_5588.n162 a_9348_5588.n161 3.229
R1394 a_9348_5588.n20 a_9348_5588.n19 3.177
R1395 a_9348_5588.n87 a_9348_5588.n86 2.984
R1396 a_9348_5588.n196 a_9348_5588.n195 2.984
R1397 a_9348_5588.n129 a_9348_5588.n126 2.87
R1398 a_9348_5588.n132 a_9348_5588.n131 2.87
R1399 a_9348_5588.n65 a_9348_5588.n64 2.87
R1400 a_9348_5588.n62 a_9348_5588.n59 2.87
R1401 a_9348_5588.n167 a_9348_5588.n165 2.87
R1402 a_9348_5588.n161 a_9348_5588.n160 2.87
R1403 a_9348_5588.n122 a_9348_5588.n121 2.511
R1404 a_9348_5588.n123 a_9348_5588.n122 2.511
R1405 a_9348_5588.n56 a_9348_5588.n55 2.511
R1406 a_9348_5588.n55 a_9348_5588.n54 2.511
R1407 a_9348_5588.n173 a_9348_5588.n170 2.511
R1408 a_9348_5588.n170 a_9348_5588.n169 2.511
R1409 a_9348_5588.n137 a_9348_5588.n134 2.152
R1410 a_9348_5588.n140 a_9348_5588.n139 2.152
R1411 a_9348_5588.n73 a_9348_5588.n72 2.152
R1412 a_9348_5588.n70 a_9348_5588.n67 2.152
R1413 a_9348_5588.n4 a_9348_5588.n1 2.152
R1414 a_9348_5588.n7 a_9348_5588.n6 2.152
R1415 a_9348_5588.n114 a_9348_5588.n113 1.794
R1416 a_9348_5588.n115 a_9348_5588.n114 1.794
R1417 a_9348_5588.n48 a_9348_5588.n47 1.794
R1418 a_9348_5588.n47 a_9348_5588.n46 1.794
R1419 a_9348_5588.n181 a_9348_5588.n178 1.794
R1420 a_9348_5588.n178 a_9348_5588.n177 1.794
R1421 a_9348_5588.n80 a_9348_5588.n77 1.076
R1422 a_9348_5588.n77 a_9348_5588.n76 1.076
R1423 a_9348_5588.n10 a_9348_5588.n9 1.076
R1424 a_9348_5588.n13 a_9348_5588.n10 1.076
R1425 a_9348_5588.n189 a_9348_5588.n186 1.076
R1426 a_9348_5588.n186 a_9348_5588.n185 1.076
R1427 a_9348_5588.n88 a_9348_5588.n85 0.358
R1428 a_9348_5588.n85 a_9348_5588.n84 0.358
R1429 a_9348_5588.n18 a_9348_5588.n17 0.358
R1430 a_9348_5588.n21 a_9348_5588.n18 0.358
R1431 a_9348_5588.n197 a_9348_5588.n194 0.358
R1432 a_9348_5588.n194 a_9348_5588.n193 0.358
R1433 a_9348_5588.n93 a_9348_5588.n92 0.144
R1434 a_9348_5588.n96 a_9348_5588.n95 0.144
R1435 a_9348_5588.n99 a_9348_5588.n98 0.144
R1436 a_9348_5588.n102 a_9348_5588.n101 0.144
R1437 a_9348_5588.n105 a_9348_5588.n104 0.144
R1438 a_9348_5588.n38 a_9348_5588.n37 0.144
R1439 a_9348_5588.n35 a_9348_5588.n34 0.144
R1440 a_9348_5588.n32 a_9348_5588.n31 0.144
R1441 a_9348_5588.n29 a_9348_5588.n28 0.144
R1442 a_9348_5588.n26 a_9348_5588.n25 0.144
R1443 a_9348_5588.n157 a_9348_5588.n156 0.144
R1444 a_9348_5588.n154 a_9348_5588.n153 0.144
R1445 a_9348_5588.n151 a_9348_5588.n150 0.144
R1446 a_9348_5588.n148 a_9348_5588.n147 0.144
R1447 a_9348_5588.n95 a_9348_5588.n94 0.038
R1448 a_9348_5588.n28 a_9348_5588.n27 0.038
R1449 a_9348_5588.n158 a_9348_5588.n157 0.038
R1450 a_9348_5588.n98 a_9348_5588.n97 0.032
R1451 a_9348_5588.n31 a_9348_5588.n30 0.032
R1452 a_9348_5588.n155 a_9348_5588.n154 0.032
R1453 a_9348_5588.n106 a_9348_5588.n105 0.029
R1454 a_9348_5588.n39 a_9348_5588.n38 0.029
R1455 a_9348_5588.n147 a_9348_5588.n146 0.029
R1456 a_9348_5588.n101 a_9348_5588.n100 0.027
R1457 a_9348_5588.n34 a_9348_5588.n33 0.027
R1458 a_9348_5588.n152 a_9348_5588.n151 0.027
R1459 a_9348_5588.n103 a_9348_5588.n102 0.024
R1460 a_9348_5588.n36 a_9348_5588.n35 0.024
R1461 a_9348_5588.n150 a_9348_5588.n149 0.024
R1462 a_9348_5588.n104 a_9348_5588.n103 0.021
R1463 a_9348_5588.n37 a_9348_5588.n36 0.021
R1464 a_9348_5588.n149 a_9348_5588.n148 0.021
R1465 a_9348_5588.n100 a_9348_5588.n99 0.019
R1466 a_9348_5588.n33 a_9348_5588.n32 0.019
R1467 a_9348_5588.n153 a_9348_5588.n152 0.019
R1468 a_9348_5588.n107 a_9348_5588.n106 0.016
R1469 a_9348_5588.n40 a_9348_5588.n39 0.016
R1470 a_9348_5588.n146 a_9348_5588.n145 0.016
R1471 a_9348_5588.n97 a_9348_5588.n96 0.013
R1472 a_9348_5588.n30 a_9348_5588.n29 0.013
R1473 a_9348_5588.n156 a_9348_5588.n155 0.013
R1474 a_9348_5588.n94 a_9348_5588.n93 0.008
R1475 a_9348_5588.n27 a_9348_5588.n26 0.008
R1476 a_9348_5588.n159 a_9348_5588.n158 0.008
R1477 a_1562_1830.n108 a_1562_1830.t5 1397.31
R1478 a_1562_1830.n118 a_1562_1830.n111 1208.44
R1479 a_1562_1830.n109 a_1562_1830.t4 1031.48
R1480 a_1562_1830.n111 a_1562_1830.n110 1031.48
R1481 a_1562_1830.n115 a_1562_1830.n114 963.661
R1482 a_1562_1830.n117 a_1562_1830.t3 948.736
R1483 a_1562_1830.n110 a_1562_1830.n107 877.239
R1484 a_1562_1830.n109 a_1562_1830.n108 877.239
R1485 a_1562_1830.n116 a_1562_1830.n112 854.746
R1486 a_1562_1830.n115 a_1562_1830.n113 841.893
R1487 a_1562_1830.n119 a_1562_1830.t2 221.859
R1488 a_1562_1830.n120 a_1562_1830.n106 186.344
R1489 a_1562_1830.n118 a_1562_1830.n117 163.738
R1490 a_1562_1830.n130 a_1562_1830.n120 163.596
R1491 a_1562_1830.n110 a_1562_1830.n109 154.24
R1492 a_1562_1830.n116 a_1562_1830.n115 137.116
R1493 a_1562_1830.n55 a_1562_1830.t1 64.755
R1494 a_1562_1830.n106 a_1562_1830.n71 49.503
R1495 a_1562_1830.t0 a_1562_1830.n130 122.225
R1496 a_1562_1830.n100 a_1562_1830.n99 32.833
R1497 a_1562_1830.t0 a_1562_1830.n39 32.727
R1498 a_1562_1830.n56 a_1562_1830.n55 30.598
R1499 a_1562_1830.n39 a_1562_1830.n1 29.09
R1500 a_1562_1830.n92 a_1562_1830.n91 26.863
R1501 a_1562_1830.n117 a_1562_1830.n116 24.1
R1502 a_1562_1830.n84 a_1562_1830.n83 20.893
R1503 a_1562_1830.n124 a_1562_1830.n123 20
R1504 a_1562_1830.n6 a_1562_1830.n5 16.363
R1505 a_1562_1830.n101 a_1562_1830.n100 15
R1506 a_1562_1830.n93 a_1562_1830.n92 15
R1507 a_1562_1830.n85 a_1562_1830.n84 15
R1508 a_1562_1830.n77 a_1562_1830.n76 15
R1509 a_1562_1830.n44 a_1562_1830.n43 15
R1510 a_1562_1830.n52 a_1562_1830.n51 15
R1511 a_1562_1830.n98 a_1562_1830.n97 15
R1512 a_1562_1830.n90 a_1562_1830.n89 15
R1513 a_1562_1830.n82 a_1562_1830.n81 15
R1514 a_1562_1830.n74 a_1562_1830.n73 15
R1515 a_1562_1830.n46 a_1562_1830.n45 15
R1516 a_1562_1830.n54 a_1562_1830.n53 15
R1517 a_1562_1830.n31 a_1562_1830.n30 15
R1518 a_1562_1830.n23 a_1562_1830.n22 15
R1519 a_1562_1830.n15 a_1562_1830.n14 15
R1520 a_1562_1830.n7 a_1562_1830.n6 15
R1521 a_1562_1830.n125 a_1562_1830.n124 15
R1522 a_1562_1830.n39 a_1562_1830.n38 15
R1523 a_1562_1830.n33 a_1562_1830.n32 15
R1524 a_1562_1830.n25 a_1562_1830.n24 15
R1525 a_1562_1830.n17 a_1562_1830.n16 15
R1526 a_1562_1830.n9 a_1562_1830.n8 15
R1527 a_1562_1830.n122 a_1562_1830.n121 15
R1528 a_1562_1830.n76 a_1562_1830.n75 14.924
R1529 a_1562_1830.n55 a_1562_1830.n54 14.123
R1530 a_1562_1830.n129 a_1562_1830.n128 13.634
R1531 a_1562_1830.n105 a_1562_1830.n104 13.544
R1532 a_1562_1830.n47 a_1562_1830.n46 12.917
R1533 a_1562_1830.n74 a_1562_1830.n72 12.917
R1534 a_1562_1830.n82 a_1562_1830.n80 12.917
R1535 a_1562_1830.n90 a_1562_1830.n88 12.917
R1536 a_1562_1830.n98 a_1562_1830.n96 12.917
R1537 a_1562_1830.n10 a_1562_1830.n9 12.917
R1538 a_1562_1830.n18 a_1562_1830.n17 12.917
R1539 a_1562_1830.n26 a_1562_1830.n25 12.917
R1540 a_1562_1830.n34 a_1562_1830.n33 12.917
R1541 a_1562_1830.n14 a_1562_1830.n13 12.727
R1542 a_1562_1830.n22 a_1562_1830.n21 9.09
R1543 a_1562_1830.n43 a_1562_1830.n42 8.954
R1544 a_1562_1830.n106 a_1562_1830.n105 8.805
R1545 a_1562_1830.n130 a_1562_1830.n129 8.695
R1546 a_1562_1830.n54 a_1562_1830.n52 5.741
R1547 a_1562_1830.n48 a_1562_1830.n47 5.741
R1548 a_1562_1830.n35 a_1562_1830.n34 5.741
R1549 a_1562_1830.n38 a_1562_1830.n37 5.741
R1550 a_1562_1830.n30 a_1562_1830.n29 5.454
R1551 a_1562_1830.n46 a_1562_1830.n44 5.023
R1552 a_1562_1830.n27 a_1562_1830.n26 5.023
R1553 a_1562_1830.n33 a_1562_1830.n31 5.023
R1554 a_1562_1830.n77 a_1562_1830.n74 4.305
R1555 a_1562_1830.n80 a_1562_1830.n79 4.305
R1556 a_1562_1830.n19 a_1562_1830.n18 4.305
R1557 a_1562_1830.n25 a_1562_1830.n23 4.305
R1558 a_1562_1830.n102 a_1562_1830.n101 3.947
R1559 a_1562_1830.n103 a_1562_1830.n102 3.947
R1560 a_1562_1830.n127 a_1562_1830.n126 3.947
R1561 a_1562_1830.n126 a_1562_1830.n125 3.947
R1562 a_1562_1830.n85 a_1562_1830.n82 3.588
R1563 a_1562_1830.n88 a_1562_1830.n87 3.588
R1564 a_1562_1830.n11 a_1562_1830.n10 3.588
R1565 a_1562_1830.n17 a_1562_1830.n15 3.588
R1566 a_1562_1830.n94 a_1562_1830.n93 3.229
R1567 a_1562_1830.n95 a_1562_1830.n94 3.229
R1568 a_1562_1830.n4 a_1562_1830.n3 3.229
R1569 a_1562_1830.n7 a_1562_1830.n4 3.229
R1570 a_1562_1830.n51 a_1562_1830.n50 2.984
R1571 a_1562_1830.n119 a_1562_1830.n118 2.875
R1572 a_1562_1830.n93 a_1562_1830.n90 2.87
R1573 a_1562_1830.n96 a_1562_1830.n95 2.87
R1574 a_1562_1830.n3 a_1562_1830.n2 2.87
R1575 a_1562_1830.n9 a_1562_1830.n7 2.87
R1576 a_1562_1830.n86 a_1562_1830.n85 2.511
R1577 a_1562_1830.n87 a_1562_1830.n86 2.511
R1578 a_1562_1830.n12 a_1562_1830.n11 2.511
R1579 a_1562_1830.n15 a_1562_1830.n12 2.511
R1580 a_1562_1830.n101 a_1562_1830.n98 2.152
R1581 a_1562_1830.n104 a_1562_1830.n103 2.152
R1582 a_1562_1830.n128 a_1562_1830.n127 2.152
R1583 a_1562_1830.n125 a_1562_1830.n122 2.152
R1584 a_1562_1830.n1 a_1562_1830.n0 1.818
R1585 a_1562_1830.n78 a_1562_1830.n77 1.794
R1586 a_1562_1830.n79 a_1562_1830.n78 1.794
R1587 a_1562_1830.n20 a_1562_1830.n19 1.794
R1588 a_1562_1830.n23 a_1562_1830.n20 1.794
R1589 a_1562_1830.n120 a_1562_1830.n119 1.149
R1590 a_1562_1830.n44 a_1562_1830.n41 1.076
R1591 a_1562_1830.n41 a_1562_1830.n40 1.076
R1592 a_1562_1830.n28 a_1562_1830.n27 1.076
R1593 a_1562_1830.n31 a_1562_1830.n28 1.076
R1594 a_1562_1830.n52 a_1562_1830.n49 0.358
R1595 a_1562_1830.n49 a_1562_1830.n48 0.358
R1596 a_1562_1830.n36 a_1562_1830.n35 0.358
R1597 a_1562_1830.n37 a_1562_1830.n36 0.358
R1598 a_1562_1830.n57 a_1562_1830.n56 0.144
R1599 a_1562_1830.n60 a_1562_1830.n59 0.144
R1600 a_1562_1830.n63 a_1562_1830.n62 0.144
R1601 a_1562_1830.n66 a_1562_1830.n65 0.144
R1602 a_1562_1830.n69 a_1562_1830.n68 0.144
R1603 a_1562_1830.n59 a_1562_1830.n58 0.038
R1604 a_1562_1830.n62 a_1562_1830.n61 0.032
R1605 a_1562_1830.n70 a_1562_1830.n69 0.029
R1606 a_1562_1830.n65 a_1562_1830.n64 0.027
R1607 a_1562_1830.n67 a_1562_1830.n66 0.024
R1608 a_1562_1830.n68 a_1562_1830.n67 0.021
R1609 a_1562_1830.n64 a_1562_1830.n63 0.019
R1610 a_1562_1830.n71 a_1562_1830.n70 0.016
R1611 a_1562_1830.n61 a_1562_1830.n60 0.013
R1612 a_1562_1830.n58 a_1562_1830.n57 0.008
R1613 a_3194_252.n174 a_3194_252.n173 346.466
R1614 a_3194_252.n184 a_3194_252.n174 312.05
R1615 a_3194_252.n174 a_3194_252.n106 165.043
R1616 a_3194_252.n106 a_3194_252.n71 49.503
R1617 a_3194_252.n173 a_3194_252.n138 49.503
R1618 a_3194_252.t1 a_3194_252.n184 122.225
R1619 a_3194_252.n122 a_3194_252.t2 44.725
R1620 a_3194_252.n55 a_3194_252.t0 44.725
R1621 a_3194_252.t1 a_3194_252.n39 32.727
R1622 a_3194_252.n123 a_3194_252.n122 29.514
R1623 a_3194_252.n56 a_3194_252.n55 29.514
R1624 a_3194_252.n39 a_3194_252.n1 29.09
R1625 a_3194_252.n100 a_3194_252.n99 21.29
R1626 a_3194_252.n167 a_3194_252.n166 21.29
R1627 a_3194_252.n178 a_3194_252.n177 20
R1628 a_3194_252.n92 a_3194_252.n91 17.419
R1629 a_3194_252.n159 a_3194_252.n158 17.419
R1630 a_3194_252.n6 a_3194_252.n5 16.363
R1631 a_3194_252.n101 a_3194_252.n100 15
R1632 a_3194_252.n93 a_3194_252.n92 15
R1633 a_3194_252.n85 a_3194_252.n84 15
R1634 a_3194_252.n77 a_3194_252.n76 15
R1635 a_3194_252.n44 a_3194_252.n43 15
R1636 a_3194_252.n52 a_3194_252.n51 15
R1637 a_3194_252.n98 a_3194_252.n97 15
R1638 a_3194_252.n90 a_3194_252.n89 15
R1639 a_3194_252.n82 a_3194_252.n81 15
R1640 a_3194_252.n74 a_3194_252.n73 15
R1641 a_3194_252.n46 a_3194_252.n45 15
R1642 a_3194_252.n54 a_3194_252.n53 15
R1643 a_3194_252.n119 a_3194_252.n118 15
R1644 a_3194_252.n111 a_3194_252.n110 15
R1645 a_3194_252.n144 a_3194_252.n143 15
R1646 a_3194_252.n152 a_3194_252.n151 15
R1647 a_3194_252.n160 a_3194_252.n159 15
R1648 a_3194_252.n168 a_3194_252.n167 15
R1649 a_3194_252.n121 a_3194_252.n120 15
R1650 a_3194_252.n113 a_3194_252.n112 15
R1651 a_3194_252.n141 a_3194_252.n140 15
R1652 a_3194_252.n149 a_3194_252.n148 15
R1653 a_3194_252.n157 a_3194_252.n156 15
R1654 a_3194_252.n165 a_3194_252.n164 15
R1655 a_3194_252.n31 a_3194_252.n30 15
R1656 a_3194_252.n23 a_3194_252.n22 15
R1657 a_3194_252.n15 a_3194_252.n14 15
R1658 a_3194_252.n7 a_3194_252.n6 15
R1659 a_3194_252.n179 a_3194_252.n178 15
R1660 a_3194_252.n39 a_3194_252.n38 15
R1661 a_3194_252.n33 a_3194_252.n32 15
R1662 a_3194_252.n25 a_3194_252.n24 15
R1663 a_3194_252.n17 a_3194_252.n16 15
R1664 a_3194_252.n9 a_3194_252.n8 15
R1665 a_3194_252.n176 a_3194_252.n175 15
R1666 a_3194_252.n55 a_3194_252.n54 14.523
R1667 a_3194_252.n122 a_3194_252.n121 14.523
R1668 a_3194_252.n183 a_3194_252.n182 13.634
R1669 a_3194_252.n105 a_3194_252.n104 13.624
R1670 a_3194_252.n172 a_3194_252.n171 13.624
R1671 a_3194_252.n84 a_3194_252.n83 13.548
R1672 a_3194_252.n151 a_3194_252.n150 13.548
R1673 a_3194_252.n47 a_3194_252.n46 12.917
R1674 a_3194_252.n74 a_3194_252.n72 12.917
R1675 a_3194_252.n82 a_3194_252.n80 12.917
R1676 a_3194_252.n90 a_3194_252.n88 12.917
R1677 a_3194_252.n98 a_3194_252.n96 12.917
R1678 a_3194_252.n165 a_3194_252.n163 12.917
R1679 a_3194_252.n157 a_3194_252.n155 12.917
R1680 a_3194_252.n149 a_3194_252.n147 12.917
R1681 a_3194_252.n141 a_3194_252.n139 12.917
R1682 a_3194_252.n114 a_3194_252.n113 12.917
R1683 a_3194_252.n10 a_3194_252.n9 12.917
R1684 a_3194_252.n18 a_3194_252.n17 12.917
R1685 a_3194_252.n26 a_3194_252.n25 12.917
R1686 a_3194_252.n34 a_3194_252.n33 12.917
R1687 a_3194_252.n14 a_3194_252.n13 12.727
R1688 a_3194_252.n76 a_3194_252.n75 9.677
R1689 a_3194_252.n143 a_3194_252.n142 9.677
R1690 a_3194_252.n22 a_3194_252.n21 9.09
R1691 a_3194_252.n106 a_3194_252.n105 8.708
R1692 a_3194_252.n173 a_3194_252.n172 8.708
R1693 a_3194_252.n184 a_3194_252.n183 8.695
R1694 a_3194_252.n43 a_3194_252.n42 5.806
R1695 a_3194_252.n110 a_3194_252.n109 5.806
R1696 a_3194_252.n54 a_3194_252.n52 5.741
R1697 a_3194_252.n48 a_3194_252.n47 5.741
R1698 a_3194_252.n115 a_3194_252.n114 5.741
R1699 a_3194_252.n121 a_3194_252.n119 5.741
R1700 a_3194_252.n35 a_3194_252.n34 5.741
R1701 a_3194_252.n38 a_3194_252.n37 5.741
R1702 a_3194_252.n30 a_3194_252.n29 5.454
R1703 a_3194_252.n46 a_3194_252.n44 5.023
R1704 a_3194_252.n113 a_3194_252.n111 5.023
R1705 a_3194_252.n27 a_3194_252.n26 5.023
R1706 a_3194_252.n33 a_3194_252.n31 5.023
R1707 a_3194_252.n77 a_3194_252.n74 4.305
R1708 a_3194_252.n80 a_3194_252.n79 4.305
R1709 a_3194_252.n147 a_3194_252.n146 4.305
R1710 a_3194_252.n144 a_3194_252.n141 4.305
R1711 a_3194_252.n19 a_3194_252.n18 4.305
R1712 a_3194_252.n25 a_3194_252.n23 4.305
R1713 a_3194_252.n102 a_3194_252.n101 3.947
R1714 a_3194_252.n103 a_3194_252.n102 3.947
R1715 a_3194_252.n170 a_3194_252.n169 3.947
R1716 a_3194_252.n169 a_3194_252.n168 3.947
R1717 a_3194_252.n181 a_3194_252.n180 3.947
R1718 a_3194_252.n180 a_3194_252.n179 3.947
R1719 a_3194_252.n85 a_3194_252.n82 3.588
R1720 a_3194_252.n88 a_3194_252.n87 3.588
R1721 a_3194_252.n155 a_3194_252.n154 3.588
R1722 a_3194_252.n152 a_3194_252.n149 3.588
R1723 a_3194_252.n11 a_3194_252.n10 3.588
R1724 a_3194_252.n17 a_3194_252.n15 3.588
R1725 a_3194_252.n94 a_3194_252.n93 3.229
R1726 a_3194_252.n95 a_3194_252.n94 3.229
R1727 a_3194_252.n162 a_3194_252.n161 3.229
R1728 a_3194_252.n161 a_3194_252.n160 3.229
R1729 a_3194_252.n4 a_3194_252.n3 3.229
R1730 a_3194_252.n7 a_3194_252.n4 3.229
R1731 a_3194_252.n93 a_3194_252.n90 2.87
R1732 a_3194_252.n96 a_3194_252.n95 2.87
R1733 a_3194_252.n163 a_3194_252.n162 2.87
R1734 a_3194_252.n160 a_3194_252.n157 2.87
R1735 a_3194_252.n3 a_3194_252.n2 2.87
R1736 a_3194_252.n9 a_3194_252.n7 2.87
R1737 a_3194_252.n86 a_3194_252.n85 2.511
R1738 a_3194_252.n87 a_3194_252.n86 2.511
R1739 a_3194_252.n154 a_3194_252.n153 2.511
R1740 a_3194_252.n153 a_3194_252.n152 2.511
R1741 a_3194_252.n12 a_3194_252.n11 2.511
R1742 a_3194_252.n15 a_3194_252.n12 2.511
R1743 a_3194_252.n101 a_3194_252.n98 2.152
R1744 a_3194_252.n104 a_3194_252.n103 2.152
R1745 a_3194_252.n171 a_3194_252.n170 2.152
R1746 a_3194_252.n168 a_3194_252.n165 2.152
R1747 a_3194_252.n182 a_3194_252.n181 2.152
R1748 a_3194_252.n179 a_3194_252.n176 2.152
R1749 a_3194_252.n51 a_3194_252.n50 1.935
R1750 a_3194_252.n118 a_3194_252.n117 1.935
R1751 a_3194_252.n1 a_3194_252.n0 1.818
R1752 a_3194_252.n78 a_3194_252.n77 1.794
R1753 a_3194_252.n79 a_3194_252.n78 1.794
R1754 a_3194_252.n146 a_3194_252.n145 1.794
R1755 a_3194_252.n145 a_3194_252.n144 1.794
R1756 a_3194_252.n20 a_3194_252.n19 1.794
R1757 a_3194_252.n23 a_3194_252.n20 1.794
R1758 a_3194_252.n44 a_3194_252.n41 1.076
R1759 a_3194_252.n41 a_3194_252.n40 1.076
R1760 a_3194_252.n108 a_3194_252.n107 1.076
R1761 a_3194_252.n111 a_3194_252.n108 1.076
R1762 a_3194_252.n28 a_3194_252.n27 1.076
R1763 a_3194_252.n31 a_3194_252.n28 1.076
R1764 a_3194_252.n52 a_3194_252.n49 0.358
R1765 a_3194_252.n49 a_3194_252.n48 0.358
R1766 a_3194_252.n116 a_3194_252.n115 0.358
R1767 a_3194_252.n119 a_3194_252.n116 0.358
R1768 a_3194_252.n36 a_3194_252.n35 0.358
R1769 a_3194_252.n37 a_3194_252.n36 0.358
R1770 a_3194_252.n57 a_3194_252.n56 0.144
R1771 a_3194_252.n60 a_3194_252.n59 0.144
R1772 a_3194_252.n63 a_3194_252.n62 0.144
R1773 a_3194_252.n66 a_3194_252.n65 0.144
R1774 a_3194_252.n69 a_3194_252.n68 0.144
R1775 a_3194_252.n136 a_3194_252.n135 0.144
R1776 a_3194_252.n133 a_3194_252.n132 0.144
R1777 a_3194_252.n130 a_3194_252.n129 0.144
R1778 a_3194_252.n127 a_3194_252.n126 0.144
R1779 a_3194_252.n124 a_3194_252.n123 0.144
R1780 a_3194_252.n59 a_3194_252.n58 0.038
R1781 a_3194_252.n126 a_3194_252.n125 0.038
R1782 a_3194_252.n62 a_3194_252.n61 0.032
R1783 a_3194_252.n129 a_3194_252.n128 0.032
R1784 a_3194_252.n70 a_3194_252.n69 0.029
R1785 a_3194_252.n137 a_3194_252.n136 0.029
R1786 a_3194_252.n65 a_3194_252.n64 0.027
R1787 a_3194_252.n132 a_3194_252.n131 0.027
R1788 a_3194_252.n67 a_3194_252.n66 0.024
R1789 a_3194_252.n134 a_3194_252.n133 0.024
R1790 a_3194_252.n68 a_3194_252.n67 0.021
R1791 a_3194_252.n135 a_3194_252.n134 0.021
R1792 a_3194_252.n64 a_3194_252.n63 0.019
R1793 a_3194_252.n131 a_3194_252.n130 0.019
R1794 a_3194_252.n71 a_3194_252.n70 0.016
R1795 a_3194_252.n138 a_3194_252.n137 0.016
R1796 a_3194_252.n61 a_3194_252.n60 0.013
R1797 a_3194_252.n128 a_3194_252.n127 0.013
R1798 a_3194_252.n58 a_3194_252.n57 0.008
R1799 a_3194_252.n125 a_3194_252.n124 0.008
R1800 a_4518_1814.n107 a_4518_1814.t5 1394.31
R1801 a_4518_1814.n118 a_4518_1814.n111 1202.83
R1802 a_4518_1814.n109 a_4518_1814.n108 1031.48
R1803 a_4518_1814.n111 a_4518_1814.n110 1031.48
R1804 a_4518_1814.n114 a_4518_1814.n113 963.661
R1805 a_4518_1814.n117 a_4518_1814.n116 948.736
R1806 a_4518_1814.n110 a_4518_1814.t3 877.239
R1807 a_4518_1814.n109 a_4518_1814.n107 877.239
R1808 a_4518_1814.n115 a_4518_1814.n112 854.746
R1809 a_4518_1814.n114 a_4518_1814.t4 841.893
R1810 a_4518_1814.n119 a_4518_1814.t0 222.024
R1811 a_4518_1814.n120 a_4518_1814.n106 186.348
R1812 a_4518_1814.n130 a_4518_1814.n120 163.592
R1813 a_4518_1814.n118 a_4518_1814.n117 162.489
R1814 a_4518_1814.n110 a_4518_1814.n109 154.24
R1815 a_4518_1814.n115 a_4518_1814.n114 137.116
R1816 a_4518_1814.n55 a_4518_1814.t2 64.755
R1817 a_4518_1814.n106 a_4518_1814.n71 49.503
R1818 a_4518_1814.t1 a_4518_1814.n130 122.225
R1819 a_4518_1814.n100 a_4518_1814.n99 32.833
R1820 a_4518_1814.t1 a_4518_1814.n39 32.727
R1821 a_4518_1814.n56 a_4518_1814.n55 30.598
R1822 a_4518_1814.n39 a_4518_1814.n1 29.09
R1823 a_4518_1814.n92 a_4518_1814.n91 26.863
R1824 a_4518_1814.n117 a_4518_1814.n115 24.1
R1825 a_4518_1814.n84 a_4518_1814.n83 20.893
R1826 a_4518_1814.n124 a_4518_1814.n123 20
R1827 a_4518_1814.n6 a_4518_1814.n5 16.363
R1828 a_4518_1814.n52 a_4518_1814.n51 15
R1829 a_4518_1814.n44 a_4518_1814.n43 15
R1830 a_4518_1814.n77 a_4518_1814.n76 15
R1831 a_4518_1814.n85 a_4518_1814.n84 15
R1832 a_4518_1814.n93 a_4518_1814.n92 15
R1833 a_4518_1814.n54 a_4518_1814.n53 15
R1834 a_4518_1814.n46 a_4518_1814.n45 15
R1835 a_4518_1814.n74 a_4518_1814.n73 15
R1836 a_4518_1814.n82 a_4518_1814.n81 15
R1837 a_4518_1814.n90 a_4518_1814.n89 15
R1838 a_4518_1814.n98 a_4518_1814.n97 15
R1839 a_4518_1814.n101 a_4518_1814.n100 15
R1840 a_4518_1814.n31 a_4518_1814.n30 15
R1841 a_4518_1814.n23 a_4518_1814.n22 15
R1842 a_4518_1814.n15 a_4518_1814.n14 15
R1843 a_4518_1814.n7 a_4518_1814.n6 15
R1844 a_4518_1814.n125 a_4518_1814.n124 15
R1845 a_4518_1814.n39 a_4518_1814.n38 15
R1846 a_4518_1814.n33 a_4518_1814.n32 15
R1847 a_4518_1814.n25 a_4518_1814.n24 15
R1848 a_4518_1814.n17 a_4518_1814.n16 15
R1849 a_4518_1814.n9 a_4518_1814.n8 15
R1850 a_4518_1814.n122 a_4518_1814.n121 15
R1851 a_4518_1814.n76 a_4518_1814.n75 14.924
R1852 a_4518_1814.n55 a_4518_1814.n54 14.123
R1853 a_4518_1814.n129 a_4518_1814.n128 13.634
R1854 a_4518_1814.n105 a_4518_1814.n104 13.544
R1855 a_4518_1814.n47 a_4518_1814.n46 12.917
R1856 a_4518_1814.n74 a_4518_1814.n72 12.917
R1857 a_4518_1814.n82 a_4518_1814.n80 12.917
R1858 a_4518_1814.n90 a_4518_1814.n88 12.917
R1859 a_4518_1814.n98 a_4518_1814.n96 12.917
R1860 a_4518_1814.n10 a_4518_1814.n9 12.917
R1861 a_4518_1814.n18 a_4518_1814.n17 12.917
R1862 a_4518_1814.n26 a_4518_1814.n25 12.917
R1863 a_4518_1814.n34 a_4518_1814.n33 12.917
R1864 a_4518_1814.n14 a_4518_1814.n13 12.727
R1865 a_4518_1814.n22 a_4518_1814.n21 9.09
R1866 a_4518_1814.n43 a_4518_1814.n42 8.954
R1867 a_4518_1814.n106 a_4518_1814.n105 8.805
R1868 a_4518_1814.n130 a_4518_1814.n129 8.695
R1869 a_4518_1814.n54 a_4518_1814.n52 5.741
R1870 a_4518_1814.n48 a_4518_1814.n47 5.741
R1871 a_4518_1814.n35 a_4518_1814.n34 5.741
R1872 a_4518_1814.n38 a_4518_1814.n37 5.741
R1873 a_4518_1814.n30 a_4518_1814.n29 5.454
R1874 a_4518_1814.n46 a_4518_1814.n44 5.023
R1875 a_4518_1814.n27 a_4518_1814.n26 5.023
R1876 a_4518_1814.n33 a_4518_1814.n31 5.023
R1877 a_4518_1814.n119 a_4518_1814.n118 4.35
R1878 a_4518_1814.n77 a_4518_1814.n74 4.305
R1879 a_4518_1814.n80 a_4518_1814.n79 4.305
R1880 a_4518_1814.n19 a_4518_1814.n18 4.305
R1881 a_4518_1814.n25 a_4518_1814.n23 4.305
R1882 a_4518_1814.n102 a_4518_1814.n101 3.947
R1883 a_4518_1814.n103 a_4518_1814.n102 3.947
R1884 a_4518_1814.n127 a_4518_1814.n126 3.947
R1885 a_4518_1814.n126 a_4518_1814.n125 3.947
R1886 a_4518_1814.n85 a_4518_1814.n82 3.588
R1887 a_4518_1814.n88 a_4518_1814.n87 3.588
R1888 a_4518_1814.n11 a_4518_1814.n10 3.588
R1889 a_4518_1814.n17 a_4518_1814.n15 3.588
R1890 a_4518_1814.n94 a_4518_1814.n93 3.229
R1891 a_4518_1814.n95 a_4518_1814.n94 3.229
R1892 a_4518_1814.n4 a_4518_1814.n3 3.229
R1893 a_4518_1814.n7 a_4518_1814.n4 3.229
R1894 a_4518_1814.n51 a_4518_1814.n50 2.984
R1895 a_4518_1814.n93 a_4518_1814.n90 2.87
R1896 a_4518_1814.n96 a_4518_1814.n95 2.87
R1897 a_4518_1814.n3 a_4518_1814.n2 2.87
R1898 a_4518_1814.n9 a_4518_1814.n7 2.87
R1899 a_4518_1814.n86 a_4518_1814.n85 2.511
R1900 a_4518_1814.n87 a_4518_1814.n86 2.511
R1901 a_4518_1814.n12 a_4518_1814.n11 2.511
R1902 a_4518_1814.n15 a_4518_1814.n12 2.511
R1903 a_4518_1814.n101 a_4518_1814.n98 2.152
R1904 a_4518_1814.n104 a_4518_1814.n103 2.152
R1905 a_4518_1814.n128 a_4518_1814.n127 2.152
R1906 a_4518_1814.n125 a_4518_1814.n122 2.152
R1907 a_4518_1814.n1 a_4518_1814.n0 1.818
R1908 a_4518_1814.n78 a_4518_1814.n77 1.794
R1909 a_4518_1814.n79 a_4518_1814.n78 1.794
R1910 a_4518_1814.n20 a_4518_1814.n19 1.794
R1911 a_4518_1814.n23 a_4518_1814.n20 1.794
R1912 a_4518_1814.n44 a_4518_1814.n41 1.076
R1913 a_4518_1814.n41 a_4518_1814.n40 1.076
R1914 a_4518_1814.n28 a_4518_1814.n27 1.076
R1915 a_4518_1814.n31 a_4518_1814.n28 1.076
R1916 a_4518_1814.n120 a_4518_1814.n119 1.036
R1917 a_4518_1814.n52 a_4518_1814.n49 0.358
R1918 a_4518_1814.n49 a_4518_1814.n48 0.358
R1919 a_4518_1814.n36 a_4518_1814.n35 0.358
R1920 a_4518_1814.n37 a_4518_1814.n36 0.358
R1921 a_4518_1814.n57 a_4518_1814.n56 0.144
R1922 a_4518_1814.n60 a_4518_1814.n59 0.144
R1923 a_4518_1814.n63 a_4518_1814.n62 0.144
R1924 a_4518_1814.n66 a_4518_1814.n65 0.144
R1925 a_4518_1814.n69 a_4518_1814.n68 0.144
R1926 a_4518_1814.n59 a_4518_1814.n58 0.038
R1927 a_4518_1814.n62 a_4518_1814.n61 0.032
R1928 a_4518_1814.n70 a_4518_1814.n69 0.029
R1929 a_4518_1814.n65 a_4518_1814.n64 0.027
R1930 a_4518_1814.n67 a_4518_1814.n66 0.024
R1931 a_4518_1814.n68 a_4518_1814.n67 0.021
R1932 a_4518_1814.n64 a_4518_1814.n63 0.019
R1933 a_4518_1814.n71 a_4518_1814.n70 0.016
R1934 a_4518_1814.n61 a_4518_1814.n60 0.013
R1935 a_4518_1814.n58 a_4518_1814.n57 0.008
R1936 VN.n141 VN.t23 1841.24
R1937 VN.n141 VN.n140 1687
R1938 VN.n282 VN.t8 1130.59
R1939 VN.n562 VN.t3 1129.87
R1940 VN.n422 VN.t10 1129.15
R1941 VN.n680 VN.t16 1128.41
R1942 VN.n138 VN.t15 1032.27
R1943 VN.t4 VN.t1 425.925
R1944 VN.t20 VN.t4 353.584
R1945 VN.n423 VN.n352 331.475
R1946 VN.n283 VN.n212 331.422
R1947 VN.n138 VN.n137 309.769
R1948 VN.n562 VN.n561 309.715
R1949 VN.n422 VN.n421 309.652
R1950 VN.t2 VN.t20 287.962
R1951 VN.n679 VN.t0 269.565
R1952 VN.n563 VN.n492 268.184
R1953 VN.n750 VN.n749 262.827
R1954 VN.t0 VN.t9 248.148
R1955 VN.n142 VN.n141 196.128
R1956 VN.n139 VN.n68 193.601
R1957 VN.n282 VN.n281 171.677
R1958 VN.n680 VN.n679 150.353
R1959 VN.n142 VN.t14 124.634
R1960 VN.t9 VN.t2 108.213
R1961 VN.n679 VN.n632 55.926
R1962 VN.n137 VN.n102 49.503
R1963 VN.n68 VN.n33 49.503
R1964 VN.n281 VN.n246 49.503
R1965 VN.n212 VN.n177 49.503
R1966 VN.n421 VN.n386 49.503
R1967 VN.n352 VN.n317 49.503
R1968 VN.n561 VN.n526 49.503
R1969 VN.n492 VN.n457 49.503
R1970 VN.n749 VN.n714 49.503
R1971 VN.n632 VN.n597 49.503
R1972 VN.t0 VN.n666 49.503
R1973 VN.n648 VN.t11 47.31
R1974 VN.n84 VN.t7 44.725
R1975 VN.n159 VN.t17 44.725
R1976 VN.n368 VN.t5 44.725
R1977 VN.n299 VN.t18 44.725
R1978 VN.n508 VN.t12 44.725
R1979 VN.n15 VN.t19 42.441
R1980 VN.n228 VN.t6 42.441
R1981 VN.n439 VN.t21 42.441
R1982 VN.n696 VN.t22 42.441
R1983 VN.n579 VN.t13 42.441
R1984 VN.n649 VN.n648 29.655
R1985 VN.n85 VN.n84 29.469
R1986 VN.n160 VN.n159 29.469
R1987 VN.n369 VN.n368 29.469
R1988 VN.n300 VN.n299 29.469
R1989 VN.n509 VN.n508 29.469
R1990 VN.n16 VN.n15 29.289
R1991 VN.n229 VN.n228 29.289
R1992 VN.n440 VN.n439 29.289
R1993 VN.n697 VN.n696 29.289
R1994 VN.n580 VN.n579 29.289
R1995 VN.n678 VN.n677 22.758
R1996 VN.n131 VN.n130 21.29
R1997 VN.n206 VN.n205 21.29
R1998 VN.n415 VN.n414 21.29
R1999 VN.n346 VN.n345 21.29
R2000 VN.n555 VN.n554 21.29
R2001 VN.n62 VN.n61 20
R2002 VN.n275 VN.n274 20
R2003 VN.n486 VN.n485 20
R2004 VN.n743 VN.n742 20
R2005 VN.n626 VN.n625 20
R2006 VN.n675 VN.n674 18.62
R2007 VN.n123 VN.n122 17.419
R2008 VN.n198 VN.n197 17.419
R2009 VN.n407 VN.n406 17.419
R2010 VN.n338 VN.n337 17.419
R2011 VN.n547 VN.n546 17.419
R2012 VN.n54 VN.n53 16.363
R2013 VN.n267 VN.n266 16.363
R2014 VN.n478 VN.n477 16.363
R2015 VN.n735 VN.n734 16.363
R2016 VN.n618 VN.n617 16.363
R2017 VN.n81 VN.n80 15
R2018 VN.n73 VN.n72 15
R2019 VN.n108 VN.n107 15
R2020 VN.n116 VN.n115 15
R2021 VN.n124 VN.n123 15
R2022 VN.n83 VN.n82 15
R2023 VN.n75 VN.n74 15
R2024 VN.n105 VN.n104 15
R2025 VN.n113 VN.n112 15
R2026 VN.n121 VN.n120 15
R2027 VN.n129 VN.n128 15
R2028 VN.n132 VN.n131 15
R2029 VN.n12 VN.n11 15
R2030 VN.n4 VN.n3 15
R2031 VN.n39 VN.n38 15
R2032 VN.n47 VN.n46 15
R2033 VN.n55 VN.n54 15
R2034 VN.n14 VN.n13 15
R2035 VN.n6 VN.n5 15
R2036 VN.n36 VN.n35 15
R2037 VN.n44 VN.n43 15
R2038 VN.n52 VN.n51 15
R2039 VN.n60 VN.n59 15
R2040 VN.n63 VN.n62 15
R2041 VN.n225 VN.n224 15
R2042 VN.n217 VN.n216 15
R2043 VN.n252 VN.n251 15
R2044 VN.n260 VN.n259 15
R2045 VN.n268 VN.n267 15
R2046 VN.n227 VN.n226 15
R2047 VN.n219 VN.n218 15
R2048 VN.n249 VN.n248 15
R2049 VN.n257 VN.n256 15
R2050 VN.n265 VN.n264 15
R2051 VN.n273 VN.n272 15
R2052 VN.n276 VN.n275 15
R2053 VN.n156 VN.n155 15
R2054 VN.n148 VN.n147 15
R2055 VN.n183 VN.n182 15
R2056 VN.n191 VN.n190 15
R2057 VN.n199 VN.n198 15
R2058 VN.n158 VN.n157 15
R2059 VN.n150 VN.n149 15
R2060 VN.n180 VN.n179 15
R2061 VN.n188 VN.n187 15
R2062 VN.n196 VN.n195 15
R2063 VN.n204 VN.n203 15
R2064 VN.n207 VN.n206 15
R2065 VN.n365 VN.n364 15
R2066 VN.n357 VN.n356 15
R2067 VN.n392 VN.n391 15
R2068 VN.n400 VN.n399 15
R2069 VN.n408 VN.n407 15
R2070 VN.n367 VN.n366 15
R2071 VN.n359 VN.n358 15
R2072 VN.n389 VN.n388 15
R2073 VN.n397 VN.n396 15
R2074 VN.n405 VN.n404 15
R2075 VN.n413 VN.n412 15
R2076 VN.n416 VN.n415 15
R2077 VN.n296 VN.n295 15
R2078 VN.n288 VN.n287 15
R2079 VN.n323 VN.n322 15
R2080 VN.n331 VN.n330 15
R2081 VN.n339 VN.n338 15
R2082 VN.n298 VN.n297 15
R2083 VN.n290 VN.n289 15
R2084 VN.n320 VN.n319 15
R2085 VN.n328 VN.n327 15
R2086 VN.n336 VN.n335 15
R2087 VN.n344 VN.n343 15
R2088 VN.n347 VN.n346 15
R2089 VN.n505 VN.n504 15
R2090 VN.n497 VN.n496 15
R2091 VN.n532 VN.n531 15
R2092 VN.n540 VN.n539 15
R2093 VN.n548 VN.n547 15
R2094 VN.n507 VN.n506 15
R2095 VN.n499 VN.n498 15
R2096 VN.n529 VN.n528 15
R2097 VN.n537 VN.n536 15
R2098 VN.n545 VN.n544 15
R2099 VN.n553 VN.n552 15
R2100 VN.n556 VN.n555 15
R2101 VN.n436 VN.n435 15
R2102 VN.n428 VN.n427 15
R2103 VN.n463 VN.n462 15
R2104 VN.n471 VN.n470 15
R2105 VN.n479 VN.n478 15
R2106 VN.n438 VN.n437 15
R2107 VN.n430 VN.n429 15
R2108 VN.n460 VN.n459 15
R2109 VN.n468 VN.n467 15
R2110 VN.n476 VN.n475 15
R2111 VN.n484 VN.n483 15
R2112 VN.n487 VN.n486 15
R2113 VN.n693 VN.n692 15
R2114 VN.n685 VN.n684 15
R2115 VN.n720 VN.n719 15
R2116 VN.n728 VN.n727 15
R2117 VN.n736 VN.n735 15
R2118 VN.n695 VN.n694 15
R2119 VN.n687 VN.n686 15
R2120 VN.n717 VN.n716 15
R2121 VN.n725 VN.n724 15
R2122 VN.n733 VN.n732 15
R2123 VN.n741 VN.n740 15
R2124 VN.n744 VN.n743 15
R2125 VN.n576 VN.n575 15
R2126 VN.n568 VN.n567 15
R2127 VN.n603 VN.n602 15
R2128 VN.n611 VN.n610 15
R2129 VN.n619 VN.n618 15
R2130 VN.n578 VN.n577 15
R2131 VN.n570 VN.n569 15
R2132 VN.n600 VN.n599 15
R2133 VN.n608 VN.n607 15
R2134 VN.n616 VN.n615 15
R2135 VN.n624 VN.n623 15
R2136 VN.n627 VN.n626 15
R2137 VN.n645 VN.n644 15
R2138 VN.n637 VN.n636 15
R2139 VN.t0 VN.n672 15
R2140 VN.t0 VN.n675 15
R2141 VN.n647 VN.n646 15
R2142 VN.n639 VN.n638 15
R2143 VN.t0 VN.n667 15
R2144 VN.t0 VN.n670 15
R2145 VN.t0 VN.n673 15
R2146 VN.t0 VN.n676 15
R2147 VN.t0 VN.n678 15
R2148 VN.t0 VN.n669 15
R2149 VN.n15 VN.n14 14.586
R2150 VN.n228 VN.n227 14.586
R2151 VN.n439 VN.n438 14.586
R2152 VN.n696 VN.n695 14.586
R2153 VN.n579 VN.n578 14.586
R2154 VN.n84 VN.n83 14.523
R2155 VN.n159 VN.n158 14.523
R2156 VN.n368 VN.n367 14.523
R2157 VN.n299 VN.n298 14.523
R2158 VN.n508 VN.n507 14.523
R2159 VN.n672 VN.n671 14.482
R2160 VN.n648 VN.n647 14.457
R2161 VN.n67 VN.n66 13.634
R2162 VN.n280 VN.n279 13.634
R2163 VN.n491 VN.n490 13.634
R2164 VN.n748 VN.n747 13.634
R2165 VN.n631 VN.n630 13.634
R2166 VN.n136 VN.n135 13.624
R2167 VN.n211 VN.n210 13.624
R2168 VN.n420 VN.n419 13.624
R2169 VN.n351 VN.n350 13.624
R2170 VN.n560 VN.n559 13.624
R2171 VN.n115 VN.n114 13.548
R2172 VN.n190 VN.n189 13.548
R2173 VN.n399 VN.n398 13.548
R2174 VN.n330 VN.n329 13.548
R2175 VN.n539 VN.n538 13.548
R2176 VN.n143 VN.n142 13.203
R2177 VN.n76 VN.n75 12.917
R2178 VN.n105 VN.n103 12.917
R2179 VN.n113 VN.n111 12.917
R2180 VN.n121 VN.n119 12.917
R2181 VN.n129 VN.n127 12.917
R2182 VN.n7 VN.n6 12.917
R2183 VN.n36 VN.n34 12.917
R2184 VN.n44 VN.n42 12.917
R2185 VN.n52 VN.n50 12.917
R2186 VN.n60 VN.n58 12.917
R2187 VN.n220 VN.n219 12.917
R2188 VN.n249 VN.n247 12.917
R2189 VN.n257 VN.n255 12.917
R2190 VN.n265 VN.n263 12.917
R2191 VN.n273 VN.n271 12.917
R2192 VN.n151 VN.n150 12.917
R2193 VN.n180 VN.n178 12.917
R2194 VN.n188 VN.n186 12.917
R2195 VN.n196 VN.n194 12.917
R2196 VN.n204 VN.n202 12.917
R2197 VN.n360 VN.n359 12.917
R2198 VN.n389 VN.n387 12.917
R2199 VN.n397 VN.n395 12.917
R2200 VN.n405 VN.n403 12.917
R2201 VN.n413 VN.n411 12.917
R2202 VN.n291 VN.n290 12.917
R2203 VN.n320 VN.n318 12.917
R2204 VN.n328 VN.n326 12.917
R2205 VN.n336 VN.n334 12.917
R2206 VN.n344 VN.n342 12.917
R2207 VN.n500 VN.n499 12.917
R2208 VN.n529 VN.n527 12.917
R2209 VN.n537 VN.n535 12.917
R2210 VN.n545 VN.n543 12.917
R2211 VN.n553 VN.n551 12.917
R2212 VN.n431 VN.n430 12.917
R2213 VN.n460 VN.n458 12.917
R2214 VN.n468 VN.n466 12.917
R2215 VN.n476 VN.n474 12.917
R2216 VN.n484 VN.n482 12.917
R2217 VN.n688 VN.n687 12.917
R2218 VN.n717 VN.n715 12.917
R2219 VN.n725 VN.n723 12.917
R2220 VN.n733 VN.n731 12.917
R2221 VN.n741 VN.n739 12.917
R2222 VN.n571 VN.n570 12.917
R2223 VN.n600 VN.n598 12.917
R2224 VN.n608 VN.n606 12.917
R2225 VN.n616 VN.n614 12.917
R2226 VN.n624 VN.n622 12.917
R2227 VN.n640 VN.n639 12.917
R2228 VN.n46 VN.n45 12.727
R2229 VN.n259 VN.n258 12.727
R2230 VN.n470 VN.n469 12.727
R2231 VN.n727 VN.n726 12.727
R2232 VN.n610 VN.n609 12.727
R2233 VN.n669 VN.n668 10.344
R2234 VN.n107 VN.n106 9.677
R2235 VN.n182 VN.n181 9.677
R2236 VN.n391 VN.n390 9.677
R2237 VN.n322 VN.n321 9.677
R2238 VN.n531 VN.n530 9.677
R2239 VN.n38 VN.n37 9.09
R2240 VN.n251 VN.n250 9.09
R2241 VN.n462 VN.n461 9.09
R2242 VN.n719 VN.n718 9.09
R2243 VN.n602 VN.n601 9.09
R2244 VN.n137 VN.n136 8.708
R2245 VN.n212 VN.n211 8.708
R2246 VN.n421 VN.n420 8.708
R2247 VN.n352 VN.n351 8.708
R2248 VN.n561 VN.n560 8.708
R2249 VN.n68 VN.n67 8.695
R2250 VN.n281 VN.n280 8.695
R2251 VN.n492 VN.n491 8.695
R2252 VN.n749 VN.n748 8.695
R2253 VN.n632 VN.n631 8.695
R2254 VN.n751 VN.n750 6.964
R2255 VN.n751 VN.n563 6.521
R2256 VN.n753 VN.n283 6.477
R2257 VN.n752 VN.n423 6.475
R2258 VN.n143 VN.n139 6.409
R2259 VN.n636 VN.n635 6.206
R2260 VN.n72 VN.n71 5.806
R2261 VN.n147 VN.n146 5.806
R2262 VN.n356 VN.n355 5.806
R2263 VN.n287 VN.n286 5.806
R2264 VN.n496 VN.n495 5.806
R2265 VN.n83 VN.n81 5.741
R2266 VN.n77 VN.n76 5.741
R2267 VN.n14 VN.n12 5.741
R2268 VN.n8 VN.n7 5.741
R2269 VN.n227 VN.n225 5.741
R2270 VN.n221 VN.n220 5.741
R2271 VN.n158 VN.n156 5.741
R2272 VN.n152 VN.n151 5.741
R2273 VN.n367 VN.n365 5.741
R2274 VN.n361 VN.n360 5.741
R2275 VN.n298 VN.n296 5.741
R2276 VN.n292 VN.n291 5.741
R2277 VN.n507 VN.n505 5.741
R2278 VN.n501 VN.n500 5.741
R2279 VN.n438 VN.n436 5.741
R2280 VN.n432 VN.n431 5.741
R2281 VN.n695 VN.n693 5.741
R2282 VN.n689 VN.n688 5.741
R2283 VN.n578 VN.n576 5.741
R2284 VN.n572 VN.n571 5.741
R2285 VN.n647 VN.n645 5.741
R2286 VN.n641 VN.n640 5.741
R2287 VN.n3 VN.n2 5.454
R2288 VN.n216 VN.n215 5.454
R2289 VN.n427 VN.n426 5.454
R2290 VN.n684 VN.n683 5.454
R2291 VN.n567 VN.n566 5.454
R2292 VN.n75 VN.n73 5.023
R2293 VN.n6 VN.n4 5.023
R2294 VN.n219 VN.n217 5.023
R2295 VN.n150 VN.n148 5.023
R2296 VN.n359 VN.n357 5.023
R2297 VN.n290 VN.n288 5.023
R2298 VN.n499 VN.n497 5.023
R2299 VN.n430 VN.n428 5.023
R2300 VN.n687 VN.n685 5.023
R2301 VN.n570 VN.n568 5.023
R2302 VN.n639 VN.n637 5.023
R2303 VN.n108 VN.n105 4.305
R2304 VN.n111 VN.n110 4.305
R2305 VN.n39 VN.n36 4.305
R2306 VN.n42 VN.n41 4.305
R2307 VN.n252 VN.n249 4.305
R2308 VN.n255 VN.n254 4.305
R2309 VN.n183 VN.n180 4.305
R2310 VN.n186 VN.n185 4.305
R2311 VN.n392 VN.n389 4.305
R2312 VN.n395 VN.n394 4.305
R2313 VN.n323 VN.n320 4.305
R2314 VN.n326 VN.n325 4.305
R2315 VN.n532 VN.n529 4.305
R2316 VN.n535 VN.n534 4.305
R2317 VN.n463 VN.n460 4.305
R2318 VN.n466 VN.n465 4.305
R2319 VN.n720 VN.n717 4.305
R2320 VN.n723 VN.n722 4.305
R2321 VN.n603 VN.n600 4.305
R2322 VN.n606 VN.n605 4.305
R2323 VN.n133 VN.n132 3.947
R2324 VN.n134 VN.n133 3.947
R2325 VN.n64 VN.n63 3.947
R2326 VN.n65 VN.n64 3.947
R2327 VN.n277 VN.n276 3.947
R2328 VN.n278 VN.n277 3.947
R2329 VN.n208 VN.n207 3.947
R2330 VN.n209 VN.n208 3.947
R2331 VN.n417 VN.n416 3.947
R2332 VN.n418 VN.n417 3.947
R2333 VN.n348 VN.n347 3.947
R2334 VN.n349 VN.n348 3.947
R2335 VN.n557 VN.n556 3.947
R2336 VN.n558 VN.n557 3.947
R2337 VN.n488 VN.n487 3.947
R2338 VN.n489 VN.n488 3.947
R2339 VN.n745 VN.n744 3.947
R2340 VN.n746 VN.n745 3.947
R2341 VN.n628 VN.n627 3.947
R2342 VN.n629 VN.n628 3.947
R2343 VN.n116 VN.n113 3.588
R2344 VN.n119 VN.n118 3.588
R2345 VN.n47 VN.n44 3.588
R2346 VN.n50 VN.n49 3.588
R2347 VN.n260 VN.n257 3.588
R2348 VN.n263 VN.n262 3.588
R2349 VN.n191 VN.n188 3.588
R2350 VN.n194 VN.n193 3.588
R2351 VN.n400 VN.n397 3.588
R2352 VN.n403 VN.n402 3.588
R2353 VN.n331 VN.n328 3.588
R2354 VN.n334 VN.n333 3.588
R2355 VN.n540 VN.n537 3.588
R2356 VN.n543 VN.n542 3.588
R2357 VN.n471 VN.n468 3.588
R2358 VN.n474 VN.n473 3.588
R2359 VN.n728 VN.n725 3.588
R2360 VN.n731 VN.n730 3.588
R2361 VN.n611 VN.n608 3.588
R2362 VN.n614 VN.n613 3.588
R2363 VN.n125 VN.n124 3.229
R2364 VN.n126 VN.n125 3.229
R2365 VN.n56 VN.n55 3.229
R2366 VN.n57 VN.n56 3.229
R2367 VN.n269 VN.n268 3.229
R2368 VN.n270 VN.n269 3.229
R2369 VN.n200 VN.n199 3.229
R2370 VN.n201 VN.n200 3.229
R2371 VN.n409 VN.n408 3.229
R2372 VN.n410 VN.n409 3.229
R2373 VN.n340 VN.n339 3.229
R2374 VN.n341 VN.n340 3.229
R2375 VN.n549 VN.n548 3.229
R2376 VN.n550 VN.n549 3.229
R2377 VN.n480 VN.n479 3.229
R2378 VN.n481 VN.n480 3.229
R2379 VN.n737 VN.n736 3.229
R2380 VN.n738 VN.n737 3.229
R2381 VN.n620 VN.n619 3.229
R2382 VN.n621 VN.n620 3.229
R2383 VN.n124 VN.n121 2.87
R2384 VN.n127 VN.n126 2.87
R2385 VN.n55 VN.n52 2.87
R2386 VN.n58 VN.n57 2.87
R2387 VN.n268 VN.n265 2.87
R2388 VN.n271 VN.n270 2.87
R2389 VN.n199 VN.n196 2.87
R2390 VN.n202 VN.n201 2.87
R2391 VN.n408 VN.n405 2.87
R2392 VN.n411 VN.n410 2.87
R2393 VN.n339 VN.n336 2.87
R2394 VN.n342 VN.n341 2.87
R2395 VN.n548 VN.n545 2.87
R2396 VN.n551 VN.n550 2.87
R2397 VN.n479 VN.n476 2.87
R2398 VN.n482 VN.n481 2.87
R2399 VN.n736 VN.n733 2.87
R2400 VN.n739 VN.n738 2.87
R2401 VN.n619 VN.n616 2.87
R2402 VN.n622 VN.n621 2.87
R2403 VN.n117 VN.n116 2.511
R2404 VN.n118 VN.n117 2.511
R2405 VN.n48 VN.n47 2.511
R2406 VN.n49 VN.n48 2.511
R2407 VN.n261 VN.n260 2.511
R2408 VN.n262 VN.n261 2.511
R2409 VN.n192 VN.n191 2.511
R2410 VN.n193 VN.n192 2.511
R2411 VN.n401 VN.n400 2.511
R2412 VN.n402 VN.n401 2.511
R2413 VN.n332 VN.n331 2.511
R2414 VN.n333 VN.n332 2.511
R2415 VN.n541 VN.n540 2.511
R2416 VN.n542 VN.n541 2.511
R2417 VN.n472 VN.n471 2.511
R2418 VN.n473 VN.n472 2.511
R2419 VN.n729 VN.n728 2.511
R2420 VN.n730 VN.n729 2.511
R2421 VN.n612 VN.n611 2.511
R2422 VN.n613 VN.n612 2.511
R2423 VN.n132 VN.n129 2.152
R2424 VN.n135 VN.n134 2.152
R2425 VN.n63 VN.n60 2.152
R2426 VN.n66 VN.n65 2.152
R2427 VN.n276 VN.n273 2.152
R2428 VN.n279 VN.n278 2.152
R2429 VN.n207 VN.n204 2.152
R2430 VN.n210 VN.n209 2.152
R2431 VN.n416 VN.n413 2.152
R2432 VN.n419 VN.n418 2.152
R2433 VN.n347 VN.n344 2.152
R2434 VN.n350 VN.n349 2.152
R2435 VN.n556 VN.n553 2.152
R2436 VN.n559 VN.n558 2.152
R2437 VN.n487 VN.n484 2.152
R2438 VN.n490 VN.n489 2.152
R2439 VN.n744 VN.n741 2.152
R2440 VN.n747 VN.n746 2.152
R2441 VN.n627 VN.n624 2.152
R2442 VN.n630 VN.n629 2.152
R2443 VN.n644 VN.n643 2.068
R2444 VN.n80 VN.n79 1.935
R2445 VN.n155 VN.n154 1.935
R2446 VN.n364 VN.n363 1.935
R2447 VN.n295 VN.n294 1.935
R2448 VN.n504 VN.n503 1.935
R2449 VN.n11 VN.n10 1.818
R2450 VN.n224 VN.n223 1.818
R2451 VN.n435 VN.n434 1.818
R2452 VN.n692 VN.n691 1.818
R2453 VN.n575 VN.n574 1.818
R2454 VN.n109 VN.n108 1.794
R2455 VN.n110 VN.n109 1.794
R2456 VN.n40 VN.n39 1.794
R2457 VN.n41 VN.n40 1.794
R2458 VN.n253 VN.n252 1.794
R2459 VN.n254 VN.n253 1.794
R2460 VN.n184 VN.n183 1.794
R2461 VN.n185 VN.n184 1.794
R2462 VN.n393 VN.n392 1.794
R2463 VN.n394 VN.n393 1.794
R2464 VN.n324 VN.n323 1.794
R2465 VN.n325 VN.n324 1.794
R2466 VN.n533 VN.n532 1.794
R2467 VN.n534 VN.n533 1.794
R2468 VN.n464 VN.n463 1.794
R2469 VN.n465 VN.n464 1.794
R2470 VN.n721 VN.n720 1.794
R2471 VN.n722 VN.n721 1.794
R2472 VN.n604 VN.n603 1.794
R2473 VN.n605 VN.n604 1.794
R2474 VN.n73 VN.n70 1.076
R2475 VN.n70 VN.n69 1.076
R2476 VN.n4 VN.n1 1.076
R2477 VN.n1 VN.n0 1.076
R2478 VN.n217 VN.n214 1.076
R2479 VN.n214 VN.n213 1.076
R2480 VN.n148 VN.n145 1.076
R2481 VN.n145 VN.n144 1.076
R2482 VN.n357 VN.n354 1.076
R2483 VN.n354 VN.n353 1.076
R2484 VN.n288 VN.n285 1.076
R2485 VN.n285 VN.n284 1.076
R2486 VN.n497 VN.n494 1.076
R2487 VN.n494 VN.n493 1.076
R2488 VN.n428 VN.n425 1.076
R2489 VN.n425 VN.n424 1.076
R2490 VN.n685 VN.n682 1.076
R2491 VN.n682 VN.n681 1.076
R2492 VN.n568 VN.n565 1.076
R2493 VN.n565 VN.n564 1.076
R2494 VN.n637 VN.n634 1.076
R2495 VN.n634 VN.n633 1.076
R2496 VN.n283 VN.n282 0.563
R2497 VN VN.n143 0.439
R2498 VN.n753 VN.n752 0.433
R2499 VN.n752 VN.n751 0.424
R2500 VN.n563 VN.n562 0.411
R2501 VN.n81 VN.n78 0.358
R2502 VN.n78 VN.n77 0.358
R2503 VN.n12 VN.n9 0.358
R2504 VN.n9 VN.n8 0.358
R2505 VN.n225 VN.n222 0.358
R2506 VN.n222 VN.n221 0.358
R2507 VN.n156 VN.n153 0.358
R2508 VN.n153 VN.n152 0.358
R2509 VN.n365 VN.n362 0.358
R2510 VN.n362 VN.n361 0.358
R2511 VN.n296 VN.n293 0.358
R2512 VN.n293 VN.n292 0.358
R2513 VN.n505 VN.n502 0.358
R2514 VN.n502 VN.n501 0.358
R2515 VN.n436 VN.n433 0.358
R2516 VN.n433 VN.n432 0.358
R2517 VN.n693 VN.n690 0.358
R2518 VN.n690 VN.n689 0.358
R2519 VN.n576 VN.n573 0.358
R2520 VN.n573 VN.n572 0.358
R2521 VN.n645 VN.n642 0.358
R2522 VN.n642 VN.n641 0.358
R2523 VN.n423 VN.n422 0.345
R2524 VN.n139 VN.n138 0.309
R2525 VN.n88 VN.n87 0.144
R2526 VN.n91 VN.n90 0.144
R2527 VN.n94 VN.n93 0.144
R2528 VN.n97 VN.n96 0.144
R2529 VN.n100 VN.n99 0.144
R2530 VN.n19 VN.n18 0.144
R2531 VN.n22 VN.n21 0.144
R2532 VN.n25 VN.n24 0.144
R2533 VN.n28 VN.n27 0.144
R2534 VN.n31 VN.n30 0.144
R2535 VN.n232 VN.n231 0.144
R2536 VN.n235 VN.n234 0.144
R2537 VN.n238 VN.n237 0.144
R2538 VN.n241 VN.n240 0.144
R2539 VN.n244 VN.n243 0.144
R2540 VN.n163 VN.n162 0.144
R2541 VN.n166 VN.n165 0.144
R2542 VN.n169 VN.n168 0.144
R2543 VN.n172 VN.n171 0.144
R2544 VN.n175 VN.n174 0.144
R2545 VN.n372 VN.n371 0.144
R2546 VN.n375 VN.n374 0.144
R2547 VN.n378 VN.n377 0.144
R2548 VN.n381 VN.n380 0.144
R2549 VN.n384 VN.n383 0.144
R2550 VN.n303 VN.n302 0.144
R2551 VN.n306 VN.n305 0.144
R2552 VN.n309 VN.n308 0.144
R2553 VN.n312 VN.n311 0.144
R2554 VN.n315 VN.n314 0.144
R2555 VN.n512 VN.n511 0.144
R2556 VN.n515 VN.n514 0.144
R2557 VN.n518 VN.n517 0.144
R2558 VN.n521 VN.n520 0.144
R2559 VN.n524 VN.n523 0.144
R2560 VN.n443 VN.n442 0.144
R2561 VN.n446 VN.n445 0.144
R2562 VN.n449 VN.n448 0.144
R2563 VN.n452 VN.n451 0.144
R2564 VN.n455 VN.n454 0.144
R2565 VN.n700 VN.n699 0.144
R2566 VN.n703 VN.n702 0.144
R2567 VN.n706 VN.n705 0.144
R2568 VN.n709 VN.n708 0.144
R2569 VN.n712 VN.n711 0.144
R2570 VN.n583 VN.n582 0.144
R2571 VN.n586 VN.n585 0.144
R2572 VN.n589 VN.n588 0.144
R2573 VN.n592 VN.n591 0.144
R2574 VN.n595 VN.n594 0.144
R2575 VN.n652 VN.n651 0.144
R2576 VN.n655 VN.n654 0.144
R2577 VN.n658 VN.n657 0.144
R2578 VN.n661 VN.n660 0.144
R2579 VN.n664 VN.n663 0.144
R2580 VN.n87 VN.n86 0.043
R2581 VN.n18 VN.n17 0.043
R2582 VN.n231 VN.n230 0.043
R2583 VN.n162 VN.n161 0.043
R2584 VN.n371 VN.n370 0.043
R2585 VN.n302 VN.n301 0.043
R2586 VN.n511 VN.n510 0.043
R2587 VN.n442 VN.n441 0.043
R2588 VN.n699 VN.n698 0.043
R2589 VN.n582 VN.n581 0.043
R2590 VN.n651 VN.n650 0.043
R2591 VN.n750 VN.n680 0.039
R2592 VN.n90 VN.n89 0.038
R2593 VN.n21 VN.n20 0.038
R2594 VN.n234 VN.n233 0.038
R2595 VN.n165 VN.n164 0.038
R2596 VN.n374 VN.n373 0.038
R2597 VN.n305 VN.n304 0.038
R2598 VN.n514 VN.n513 0.038
R2599 VN.n445 VN.n444 0.038
R2600 VN.n702 VN.n701 0.038
R2601 VN.n585 VN.n584 0.038
R2602 VN.n654 VN.n653 0.038
R2603 VN.n93 VN.n92 0.032
R2604 VN.n24 VN.n23 0.032
R2605 VN.n237 VN.n236 0.032
R2606 VN.n168 VN.n167 0.032
R2607 VN.n377 VN.n376 0.032
R2608 VN.n308 VN.n307 0.032
R2609 VN.n517 VN.n516 0.032
R2610 VN.n448 VN.n447 0.032
R2611 VN.n705 VN.n704 0.032
R2612 VN.n588 VN.n587 0.032
R2613 VN.n657 VN.n656 0.032
R2614 VN.n101 VN.n100 0.029
R2615 VN.n32 VN.n31 0.029
R2616 VN.n245 VN.n244 0.029
R2617 VN.n176 VN.n175 0.029
R2618 VN.n385 VN.n384 0.029
R2619 VN.n316 VN.n315 0.029
R2620 VN.n525 VN.n524 0.029
R2621 VN.n456 VN.n455 0.029
R2622 VN.n713 VN.n712 0.029
R2623 VN.n596 VN.n595 0.029
R2624 VN.n665 VN.n664 0.029
R2625 VN.n96 VN.n95 0.027
R2626 VN.n27 VN.n26 0.027
R2627 VN.n240 VN.n239 0.027
R2628 VN.n171 VN.n170 0.027
R2629 VN.n380 VN.n379 0.027
R2630 VN.n311 VN.n310 0.027
R2631 VN.n520 VN.n519 0.027
R2632 VN.n451 VN.n450 0.027
R2633 VN.n708 VN.n707 0.027
R2634 VN.n591 VN.n590 0.027
R2635 VN.n660 VN.n659 0.027
R2636 VN.n98 VN.n97 0.024
R2637 VN.n29 VN.n28 0.024
R2638 VN.n242 VN.n241 0.024
R2639 VN.n173 VN.n172 0.024
R2640 VN.n382 VN.n381 0.024
R2641 VN.n313 VN.n312 0.024
R2642 VN.n522 VN.n521 0.024
R2643 VN.n453 VN.n452 0.024
R2644 VN.n710 VN.n709 0.024
R2645 VN.n593 VN.n592 0.024
R2646 VN.n662 VN.n661 0.024
R2647 VN.n99 VN.n98 0.021
R2648 VN.n30 VN.n29 0.021
R2649 VN.n243 VN.n242 0.021
R2650 VN.n174 VN.n173 0.021
R2651 VN.n383 VN.n382 0.021
R2652 VN.n314 VN.n313 0.021
R2653 VN.n523 VN.n522 0.021
R2654 VN.n454 VN.n453 0.021
R2655 VN.n711 VN.n710 0.021
R2656 VN.n594 VN.n593 0.021
R2657 VN.n663 VN.n662 0.021
R2658 VN.n95 VN.n94 0.019
R2659 VN.n26 VN.n25 0.019
R2660 VN.n239 VN.n238 0.019
R2661 VN.n170 VN.n169 0.019
R2662 VN.n379 VN.n378 0.019
R2663 VN.n310 VN.n309 0.019
R2664 VN.n519 VN.n518 0.019
R2665 VN.n450 VN.n449 0.019
R2666 VN.n707 VN.n706 0.019
R2667 VN.n590 VN.n589 0.019
R2668 VN.n659 VN.n658 0.019
R2669 VN VN.n753 0.018
R2670 VN.n102 VN.n101 0.016
R2671 VN.n33 VN.n32 0.016
R2672 VN.n246 VN.n245 0.016
R2673 VN.n177 VN.n176 0.016
R2674 VN.n386 VN.n385 0.016
R2675 VN.n317 VN.n316 0.016
R2676 VN.n526 VN.n525 0.016
R2677 VN.n457 VN.n456 0.016
R2678 VN.n714 VN.n713 0.016
R2679 VN.n597 VN.n596 0.016
R2680 VN.n666 VN.n665 0.016
R2681 VN.n92 VN.n91 0.013
R2682 VN.n23 VN.n22 0.013
R2683 VN.n236 VN.n235 0.013
R2684 VN.n167 VN.n166 0.013
R2685 VN.n376 VN.n375 0.013
R2686 VN.n307 VN.n306 0.013
R2687 VN.n516 VN.n515 0.013
R2688 VN.n447 VN.n446 0.013
R2689 VN.n704 VN.n703 0.013
R2690 VN.n587 VN.n586 0.013
R2691 VN.n656 VN.n655 0.013
R2692 VN.n89 VN.n88 0.008
R2693 VN.n20 VN.n19 0.008
R2694 VN.n233 VN.n232 0.008
R2695 VN.n164 VN.n163 0.008
R2696 VN.n373 VN.n372 0.008
R2697 VN.n304 VN.n303 0.008
R2698 VN.n513 VN.n512 0.008
R2699 VN.n444 VN.n443 0.008
R2700 VN.n701 VN.n700 0.008
R2701 VN.n584 VN.n583 0.008
R2702 VN.n653 VN.n652 0.008
R2703 VN.n86 VN.n85 0.002
R2704 VN.n17 VN.n16 0.002
R2705 VN.n230 VN.n229 0.002
R2706 VN.n161 VN.n160 0.002
R2707 VN.n370 VN.n369 0.002
R2708 VN.n301 VN.n300 0.002
R2709 VN.n510 VN.n509 0.002
R2710 VN.n441 VN.n440 0.002
R2711 VN.n698 VN.n697 0.002
R2712 VN.n581 VN.n580 0.002
R2713 VN.n650 VN.n649 0.002
R2714 a_274_5606.n144 a_274_5606.n143 298.331
R2715 a_274_5606.n143 a_274_5606.n142 187.172
R2716 a_274_5606.n143 a_274_5606.n75 169.436
R2717 a_274_5606.n24 a_274_5606.t2 68.375
R2718 a_274_5606.n91 a_274_5606.t1 64.755
R2719 a_274_5606.t0 a_274_5606.n199 53.727
R2720 a_274_5606.n142 a_274_5606.n107 49.503
R2721 a_274_5606.n75 a_274_5606.n40 49.503
R2722 a_274_5606.n145 a_274_5606.n144 49.503
R2723 a_274_5606.n69 a_274_5606.n68 34.951
R2724 a_274_5606.n136 a_274_5606.n135 32.833
R2725 a_274_5606.n3 a_274_5606.n2 32.833
R2726 a_274_5606.n25 a_274_5606.n24 30.732
R2727 a_274_5606.n92 a_274_5606.n91 30.598
R2728 a_274_5606.t0 a_274_5606.n159 95.496
R2729 a_274_5606.n61 a_274_5606.n60 28.596
R2730 a_274_5606.n128 a_274_5606.n127 26.863
R2731 a_274_5606.n164 a_274_5606.n163 26.863
R2732 a_274_5606.n53 a_274_5606.n52 22.241
R2733 a_274_5606.n120 a_274_5606.n119 20.893
R2734 a_274_5606.n172 a_274_5606.n171 20.893
R2735 a_274_5606.n45 a_274_5606.n44 15.887
R2736 a_274_5606.n88 a_274_5606.n87 15
R2737 a_274_5606.n80 a_274_5606.n79 15
R2738 a_274_5606.n113 a_274_5606.n112 15
R2739 a_274_5606.n121 a_274_5606.n120 15
R2740 a_274_5606.n129 a_274_5606.n128 15
R2741 a_274_5606.n90 a_274_5606.n89 15
R2742 a_274_5606.n82 a_274_5606.n81 15
R2743 a_274_5606.n110 a_274_5606.n109 15
R2744 a_274_5606.n118 a_274_5606.n117 15
R2745 a_274_5606.n126 a_274_5606.n125 15
R2746 a_274_5606.n134 a_274_5606.n133 15
R2747 a_274_5606.n137 a_274_5606.n136 15
R2748 a_274_5606.n21 a_274_5606.n20 15
R2749 a_274_5606.n13 a_274_5606.n12 15
R2750 a_274_5606.n46 a_274_5606.n45 15
R2751 a_274_5606.n54 a_274_5606.n53 15
R2752 a_274_5606.n62 a_274_5606.n61 15
R2753 a_274_5606.n70 a_274_5606.n69 15
R2754 a_274_5606.n23 a_274_5606.n22 15
R2755 a_274_5606.n15 a_274_5606.n14 15
R2756 a_274_5606.n43 a_274_5606.n42 15
R2757 a_274_5606.n51 a_274_5606.n50 15
R2758 a_274_5606.n59 a_274_5606.n58 15
R2759 a_274_5606.n67 a_274_5606.n66 15
R2760 a_274_5606.n197 a_274_5606.n196 15
R2761 a_274_5606.n189 a_274_5606.n188 15
R2762 a_274_5606.n181 a_274_5606.n180 15
R2763 a_274_5606.n173 a_274_5606.n172 15
R2764 a_274_5606.n165 a_274_5606.n164 15
R2765 a_274_5606.n199 a_274_5606.n198 15
R2766 a_274_5606.n191 a_274_5606.n190 15
R2767 a_274_5606.n183 a_274_5606.n182 15
R2768 a_274_5606.n175 a_274_5606.n174 15
R2769 a_274_5606.n167 a_274_5606.n166 15
R2770 a_274_5606.n1 a_274_5606.n0 15
R2771 a_274_5606.n4 a_274_5606.n3 15
R2772 a_274_5606.n112 a_274_5606.n111 14.924
R2773 a_274_5606.n180 a_274_5606.n179 14.924
R2774 a_274_5606.n91 a_274_5606.n90 14.123
R2775 a_274_5606.n24 a_274_5606.n23 14.071
R2776 a_274_5606.n141 a_274_5606.n140 13.544
R2777 a_274_5606.n8 a_274_5606.n7 13.544
R2778 a_274_5606.n74 a_274_5606.n73 13.532
R2779 a_274_5606.n83 a_274_5606.n82 12.917
R2780 a_274_5606.n110 a_274_5606.n108 12.917
R2781 a_274_5606.n118 a_274_5606.n116 12.917
R2782 a_274_5606.n126 a_274_5606.n124 12.917
R2783 a_274_5606.n134 a_274_5606.n132 12.917
R2784 a_274_5606.n67 a_274_5606.n65 12.917
R2785 a_274_5606.n59 a_274_5606.n57 12.917
R2786 a_274_5606.n51 a_274_5606.n49 12.917
R2787 a_274_5606.n43 a_274_5606.n41 12.917
R2788 a_274_5606.n16 a_274_5606.n15 12.917
R2789 a_274_5606.n192 a_274_5606.n191 12.917
R2790 a_274_5606.n184 a_274_5606.n183 12.917
R2791 a_274_5606.n176 a_274_5606.n175 12.917
R2792 a_274_5606.n168 a_274_5606.n167 12.917
R2793 a_274_5606.n12 a_274_5606.n11 9.532
R2794 a_274_5606.n79 a_274_5606.n78 8.954
R2795 a_274_5606.n188 a_274_5606.n187 8.954
R2796 a_274_5606.n75 a_274_5606.n74 8.82
R2797 a_274_5606.n142 a_274_5606.n141 8.805
R2798 a_274_5606.n144 a_274_5606.n8 8.805
R2799 a_274_5606.n90 a_274_5606.n88 5.741
R2800 a_274_5606.n84 a_274_5606.n83 5.741
R2801 a_274_5606.n17 a_274_5606.n16 5.741
R2802 a_274_5606.n23 a_274_5606.n21 5.741
R2803 a_274_5606.n198 a_274_5606.n197 5.741
R2804 a_274_5606.n193 a_274_5606.n192 5.741
R2805 a_274_5606.n82 a_274_5606.n80 5.023
R2806 a_274_5606.n15 a_274_5606.n13 5.023
R2807 a_274_5606.n191 a_274_5606.n189 5.023
R2808 a_274_5606.n185 a_274_5606.n184 5.023
R2809 a_274_5606.n113 a_274_5606.n110 4.305
R2810 a_274_5606.n116 a_274_5606.n115 4.305
R2811 a_274_5606.n49 a_274_5606.n48 4.305
R2812 a_274_5606.n46 a_274_5606.n43 4.305
R2813 a_274_5606.n183 a_274_5606.n181 4.305
R2814 a_274_5606.n177 a_274_5606.n176 4.305
R2815 a_274_5606.n138 a_274_5606.n137 3.947
R2816 a_274_5606.n139 a_274_5606.n138 3.947
R2817 a_274_5606.n72 a_274_5606.n71 3.947
R2818 a_274_5606.n71 a_274_5606.n70 3.947
R2819 a_274_5606.n5 a_274_5606.n4 3.947
R2820 a_274_5606.n6 a_274_5606.n5 3.947
R2821 a_274_5606.n121 a_274_5606.n118 3.588
R2822 a_274_5606.n124 a_274_5606.n123 3.588
R2823 a_274_5606.n57 a_274_5606.n56 3.588
R2824 a_274_5606.n54 a_274_5606.n51 3.588
R2825 a_274_5606.n175 a_274_5606.n173 3.588
R2826 a_274_5606.n169 a_274_5606.n168 3.588
R2827 a_274_5606.n130 a_274_5606.n129 3.229
R2828 a_274_5606.n131 a_274_5606.n130 3.229
R2829 a_274_5606.n64 a_274_5606.n63 3.229
R2830 a_274_5606.n63 a_274_5606.n62 3.229
R2831 a_274_5606.n165 a_274_5606.n162 3.229
R2832 a_274_5606.n162 a_274_5606.n161 3.229
R2833 a_274_5606.n20 a_274_5606.n19 3.177
R2834 a_274_5606.n87 a_274_5606.n86 2.984
R2835 a_274_5606.n196 a_274_5606.n195 2.984
R2836 a_274_5606.n129 a_274_5606.n126 2.87
R2837 a_274_5606.n132 a_274_5606.n131 2.87
R2838 a_274_5606.n65 a_274_5606.n64 2.87
R2839 a_274_5606.n62 a_274_5606.n59 2.87
R2840 a_274_5606.n167 a_274_5606.n165 2.87
R2841 a_274_5606.n161 a_274_5606.n160 2.87
R2842 a_274_5606.n122 a_274_5606.n121 2.511
R2843 a_274_5606.n123 a_274_5606.n122 2.511
R2844 a_274_5606.n56 a_274_5606.n55 2.511
R2845 a_274_5606.n55 a_274_5606.n54 2.511
R2846 a_274_5606.n173 a_274_5606.n170 2.511
R2847 a_274_5606.n170 a_274_5606.n169 2.511
R2848 a_274_5606.n137 a_274_5606.n134 2.152
R2849 a_274_5606.n140 a_274_5606.n139 2.152
R2850 a_274_5606.n73 a_274_5606.n72 2.152
R2851 a_274_5606.n70 a_274_5606.n67 2.152
R2852 a_274_5606.n4 a_274_5606.n1 2.152
R2853 a_274_5606.n7 a_274_5606.n6 2.152
R2854 a_274_5606.n114 a_274_5606.n113 1.794
R2855 a_274_5606.n115 a_274_5606.n114 1.794
R2856 a_274_5606.n48 a_274_5606.n47 1.794
R2857 a_274_5606.n47 a_274_5606.n46 1.794
R2858 a_274_5606.n181 a_274_5606.n178 1.794
R2859 a_274_5606.n178 a_274_5606.n177 1.794
R2860 a_274_5606.n80 a_274_5606.n77 1.076
R2861 a_274_5606.n77 a_274_5606.n76 1.076
R2862 a_274_5606.n10 a_274_5606.n9 1.076
R2863 a_274_5606.n13 a_274_5606.n10 1.076
R2864 a_274_5606.n189 a_274_5606.n186 1.076
R2865 a_274_5606.n186 a_274_5606.n185 1.076
R2866 a_274_5606.n88 a_274_5606.n85 0.358
R2867 a_274_5606.n85 a_274_5606.n84 0.358
R2868 a_274_5606.n18 a_274_5606.n17 0.358
R2869 a_274_5606.n21 a_274_5606.n18 0.358
R2870 a_274_5606.n197 a_274_5606.n194 0.358
R2871 a_274_5606.n194 a_274_5606.n193 0.358
R2872 a_274_5606.n93 a_274_5606.n92 0.144
R2873 a_274_5606.n96 a_274_5606.n95 0.144
R2874 a_274_5606.n99 a_274_5606.n98 0.144
R2875 a_274_5606.n102 a_274_5606.n101 0.144
R2876 a_274_5606.n105 a_274_5606.n104 0.144
R2877 a_274_5606.n38 a_274_5606.n37 0.144
R2878 a_274_5606.n35 a_274_5606.n34 0.144
R2879 a_274_5606.n32 a_274_5606.n31 0.144
R2880 a_274_5606.n29 a_274_5606.n28 0.144
R2881 a_274_5606.n26 a_274_5606.n25 0.144
R2882 a_274_5606.n157 a_274_5606.n156 0.144
R2883 a_274_5606.n154 a_274_5606.n153 0.144
R2884 a_274_5606.n151 a_274_5606.n150 0.144
R2885 a_274_5606.n148 a_274_5606.n147 0.144
R2886 a_274_5606.n95 a_274_5606.n94 0.038
R2887 a_274_5606.n28 a_274_5606.n27 0.038
R2888 a_274_5606.n158 a_274_5606.n157 0.038
R2889 a_274_5606.n98 a_274_5606.n97 0.032
R2890 a_274_5606.n31 a_274_5606.n30 0.032
R2891 a_274_5606.n155 a_274_5606.n154 0.032
R2892 a_274_5606.n106 a_274_5606.n105 0.029
R2893 a_274_5606.n39 a_274_5606.n38 0.029
R2894 a_274_5606.n147 a_274_5606.n146 0.029
R2895 a_274_5606.n101 a_274_5606.n100 0.027
R2896 a_274_5606.n34 a_274_5606.n33 0.027
R2897 a_274_5606.n152 a_274_5606.n151 0.027
R2898 a_274_5606.n103 a_274_5606.n102 0.024
R2899 a_274_5606.n36 a_274_5606.n35 0.024
R2900 a_274_5606.n150 a_274_5606.n149 0.024
R2901 a_274_5606.n104 a_274_5606.n103 0.021
R2902 a_274_5606.n37 a_274_5606.n36 0.021
R2903 a_274_5606.n149 a_274_5606.n148 0.021
R2904 a_274_5606.n100 a_274_5606.n99 0.019
R2905 a_274_5606.n33 a_274_5606.n32 0.019
R2906 a_274_5606.n153 a_274_5606.n152 0.019
R2907 a_274_5606.n107 a_274_5606.n106 0.016
R2908 a_274_5606.n40 a_274_5606.n39 0.016
R2909 a_274_5606.n146 a_274_5606.n145 0.016
R2910 a_274_5606.n97 a_274_5606.n96 0.013
R2911 a_274_5606.n30 a_274_5606.n29 0.013
R2912 a_274_5606.n156 a_274_5606.n155 0.013
R2913 a_274_5606.n94 a_274_5606.n93 0.008
R2914 a_274_5606.n27 a_274_5606.n26 0.008
R2915 a_274_5606.n159 a_274_5606.n158 0.008
R2916 a_1534_3844.n112 a_1534_3844.n111 1193.37
R2917 a_1534_3844.n109 a_1534_3844.t4 1031.48
R2918 a_1534_3844.n110 a_1534_3844.n107 1031.48
R2919 a_1534_3844.n117 a_1534_3844.n116 963.661
R2920 a_1534_3844.n119 a_1534_3844.t3 948.736
R2921 a_1534_3844.n109 a_1534_3844.n108 877.239
R2922 a_1534_3844.n111 a_1534_3844.n110 877.239
R2923 a_1534_3844.n118 a_1534_3844.n114 854.746
R2924 a_1534_3844.n117 a_1534_3844.n115 841.893
R2925 a_1534_3844.n120 a_1534_3844.t0 221.783
R2926 a_1534_3844.n112 a_1534_3844.t5 207.728
R2927 a_1534_3844.n113 a_1534_3844.n106 185.413
R2928 a_1534_3844.n120 a_1534_3844.n119 166.745
R2929 a_1534_3844.n131 a_1534_3844.n121 163.552
R2930 a_1534_3844.n110 a_1534_3844.n109 154.24
R2931 a_1534_3844.n118 a_1534_3844.n117 137.116
R2932 a_1534_3844.n55 a_1534_3844.t1 64.755
R2933 a_1534_3844.n106 a_1534_3844.n71 49.503
R2934 a_1534_3844.t2 a_1534_3844.n131 122.225
R2935 a_1534_3844.n100 a_1534_3844.n99 32.833
R2936 a_1534_3844.t2 a_1534_3844.n39 32.727
R2937 a_1534_3844.n56 a_1534_3844.n55 30.598
R2938 a_1534_3844.n39 a_1534_3844.n1 29.09
R2939 a_1534_3844.n92 a_1534_3844.n91 26.863
R2940 a_1534_3844.n119 a_1534_3844.n118 24.1
R2941 a_1534_3844.n84 a_1534_3844.n83 20.893
R2942 a_1534_3844.n125 a_1534_3844.n124 20
R2943 a_1534_3844.n6 a_1534_3844.n5 16.363
R2944 a_1534_3844.n52 a_1534_3844.n51 15
R2945 a_1534_3844.n44 a_1534_3844.n43 15
R2946 a_1534_3844.n77 a_1534_3844.n76 15
R2947 a_1534_3844.n85 a_1534_3844.n84 15
R2948 a_1534_3844.n93 a_1534_3844.n92 15
R2949 a_1534_3844.n54 a_1534_3844.n53 15
R2950 a_1534_3844.n46 a_1534_3844.n45 15
R2951 a_1534_3844.n74 a_1534_3844.n73 15
R2952 a_1534_3844.n82 a_1534_3844.n81 15
R2953 a_1534_3844.n90 a_1534_3844.n89 15
R2954 a_1534_3844.n98 a_1534_3844.n97 15
R2955 a_1534_3844.n101 a_1534_3844.n100 15
R2956 a_1534_3844.n31 a_1534_3844.n30 15
R2957 a_1534_3844.n23 a_1534_3844.n22 15
R2958 a_1534_3844.n15 a_1534_3844.n14 15
R2959 a_1534_3844.n7 a_1534_3844.n6 15
R2960 a_1534_3844.n126 a_1534_3844.n125 15
R2961 a_1534_3844.n39 a_1534_3844.n38 15
R2962 a_1534_3844.n33 a_1534_3844.n32 15
R2963 a_1534_3844.n25 a_1534_3844.n24 15
R2964 a_1534_3844.n17 a_1534_3844.n16 15
R2965 a_1534_3844.n9 a_1534_3844.n8 15
R2966 a_1534_3844.n123 a_1534_3844.n122 15
R2967 a_1534_3844.n76 a_1534_3844.n75 14.924
R2968 a_1534_3844.n55 a_1534_3844.n54 14.123
R2969 a_1534_3844.n130 a_1534_3844.n129 13.634
R2970 a_1534_3844.n105 a_1534_3844.n104 13.544
R2971 a_1534_3844.n47 a_1534_3844.n46 12.917
R2972 a_1534_3844.n74 a_1534_3844.n72 12.917
R2973 a_1534_3844.n82 a_1534_3844.n80 12.917
R2974 a_1534_3844.n90 a_1534_3844.n88 12.917
R2975 a_1534_3844.n98 a_1534_3844.n96 12.917
R2976 a_1534_3844.n10 a_1534_3844.n9 12.917
R2977 a_1534_3844.n18 a_1534_3844.n17 12.917
R2978 a_1534_3844.n26 a_1534_3844.n25 12.917
R2979 a_1534_3844.n34 a_1534_3844.n33 12.917
R2980 a_1534_3844.n14 a_1534_3844.n13 12.727
R2981 a_1534_3844.n113 a_1534_3844.n112 12.141
R2982 a_1534_3844.n22 a_1534_3844.n21 9.09
R2983 a_1534_3844.n43 a_1534_3844.n42 8.954
R2984 a_1534_3844.n106 a_1534_3844.n105 8.805
R2985 a_1534_3844.n131 a_1534_3844.n130 8.695
R2986 a_1534_3844.n54 a_1534_3844.n52 5.741
R2987 a_1534_3844.n48 a_1534_3844.n47 5.741
R2988 a_1534_3844.n35 a_1534_3844.n34 5.741
R2989 a_1534_3844.n38 a_1534_3844.n37 5.741
R2990 a_1534_3844.n30 a_1534_3844.n29 5.454
R2991 a_1534_3844.n46 a_1534_3844.n44 5.023
R2992 a_1534_3844.n27 a_1534_3844.n26 5.023
R2993 a_1534_3844.n33 a_1534_3844.n31 5.023
R2994 a_1534_3844.n77 a_1534_3844.n74 4.305
R2995 a_1534_3844.n80 a_1534_3844.n79 4.305
R2996 a_1534_3844.n19 a_1534_3844.n18 4.305
R2997 a_1534_3844.n25 a_1534_3844.n23 4.305
R2998 a_1534_3844.n102 a_1534_3844.n101 3.947
R2999 a_1534_3844.n103 a_1534_3844.n102 3.947
R3000 a_1534_3844.n128 a_1534_3844.n127 3.947
R3001 a_1534_3844.n127 a_1534_3844.n126 3.947
R3002 a_1534_3844.n85 a_1534_3844.n82 3.588
R3003 a_1534_3844.n88 a_1534_3844.n87 3.588
R3004 a_1534_3844.n11 a_1534_3844.n10 3.588
R3005 a_1534_3844.n17 a_1534_3844.n15 3.588
R3006 a_1534_3844.n94 a_1534_3844.n93 3.229
R3007 a_1534_3844.n95 a_1534_3844.n94 3.229
R3008 a_1534_3844.n4 a_1534_3844.n3 3.229
R3009 a_1534_3844.n7 a_1534_3844.n4 3.229
R3010 a_1534_3844.n51 a_1534_3844.n50 2.984
R3011 a_1534_3844.n93 a_1534_3844.n90 2.87
R3012 a_1534_3844.n96 a_1534_3844.n95 2.87
R3013 a_1534_3844.n3 a_1534_3844.n2 2.87
R3014 a_1534_3844.n9 a_1534_3844.n7 2.87
R3015 a_1534_3844.n86 a_1534_3844.n85 2.511
R3016 a_1534_3844.n87 a_1534_3844.n86 2.511
R3017 a_1534_3844.n12 a_1534_3844.n11 2.511
R3018 a_1534_3844.n15 a_1534_3844.n12 2.511
R3019 a_1534_3844.n101 a_1534_3844.n98 2.152
R3020 a_1534_3844.n104 a_1534_3844.n103 2.152
R3021 a_1534_3844.n129 a_1534_3844.n128 2.152
R3022 a_1534_3844.n126 a_1534_3844.n123 2.152
R3023 a_1534_3844.n1 a_1534_3844.n0 1.818
R3024 a_1534_3844.n78 a_1534_3844.n77 1.794
R3025 a_1534_3844.n79 a_1534_3844.n78 1.794
R3026 a_1534_3844.n20 a_1534_3844.n19 1.794
R3027 a_1534_3844.n23 a_1534_3844.n20 1.794
R3028 a_1534_3844.n121 a_1534_3844.n120 1.177
R3029 a_1534_3844.n44 a_1534_3844.n41 1.076
R3030 a_1534_3844.n41 a_1534_3844.n40 1.076
R3031 a_1534_3844.n28 a_1534_3844.n27 1.076
R3032 a_1534_3844.n31 a_1534_3844.n28 1.076
R3033 a_1534_3844.n121 a_1534_3844.n113 0.85
R3034 a_1534_3844.n52 a_1534_3844.n49 0.358
R3035 a_1534_3844.n49 a_1534_3844.n48 0.358
R3036 a_1534_3844.n36 a_1534_3844.n35 0.358
R3037 a_1534_3844.n37 a_1534_3844.n36 0.358
R3038 a_1534_3844.n57 a_1534_3844.n56 0.144
R3039 a_1534_3844.n60 a_1534_3844.n59 0.144
R3040 a_1534_3844.n63 a_1534_3844.n62 0.144
R3041 a_1534_3844.n66 a_1534_3844.n65 0.144
R3042 a_1534_3844.n69 a_1534_3844.n68 0.144
R3043 a_1534_3844.n59 a_1534_3844.n58 0.038
R3044 a_1534_3844.n62 a_1534_3844.n61 0.032
R3045 a_1534_3844.n70 a_1534_3844.n69 0.029
R3046 a_1534_3844.n65 a_1534_3844.n64 0.027
R3047 a_1534_3844.n67 a_1534_3844.n66 0.024
R3048 a_1534_3844.n68 a_1534_3844.n67 0.021
R3049 a_1534_3844.n64 a_1534_3844.n63 0.019
R3050 a_1534_3844.n71 a_1534_3844.n70 0.016
R3051 a_1534_3844.n61 a_1534_3844.n60 0.013
R3052 a_1534_3844.n58 a_1534_3844.n57 0.008
R3053 a_9312_250.n174 a_9312_250.n173 273.235
R3054 a_9312_250.n184 a_9312_250.n174 243.12
R3055 a_9312_250.n174 a_9312_250.n106 165.043
R3056 a_9312_250.n106 a_9312_250.n71 49.503
R3057 a_9312_250.n173 a_9312_250.n138 49.503
R3058 a_9312_250.t0 a_9312_250.n184 122.225
R3059 a_9312_250.n55 a_9312_250.t1 44.725
R3060 a_9312_250.n122 a_9312_250.t2 42.441
R3061 a_9312_250.t0 a_9312_250.n39 32.727
R3062 a_9312_250.n56 a_9312_250.n55 29.514
R3063 a_9312_250.n123 a_9312_250.n122 29.334
R3064 a_9312_250.n39 a_9312_250.n1 29.09
R3065 a_9312_250.n100 a_9312_250.n99 21.29
R3066 a_9312_250.n167 a_9312_250.n166 20
R3067 a_9312_250.n178 a_9312_250.n177 20
R3068 a_9312_250.n92 a_9312_250.n91 17.419
R3069 a_9312_250.n159 a_9312_250.n158 16.363
R3070 a_9312_250.n6 a_9312_250.n5 16.363
R3071 a_9312_250.n101 a_9312_250.n100 15
R3072 a_9312_250.n93 a_9312_250.n92 15
R3073 a_9312_250.n85 a_9312_250.n84 15
R3074 a_9312_250.n77 a_9312_250.n76 15
R3075 a_9312_250.n44 a_9312_250.n43 15
R3076 a_9312_250.n52 a_9312_250.n51 15
R3077 a_9312_250.n98 a_9312_250.n97 15
R3078 a_9312_250.n90 a_9312_250.n89 15
R3079 a_9312_250.n82 a_9312_250.n81 15
R3080 a_9312_250.n74 a_9312_250.n73 15
R3081 a_9312_250.n46 a_9312_250.n45 15
R3082 a_9312_250.n54 a_9312_250.n53 15
R3083 a_9312_250.n119 a_9312_250.n118 15
R3084 a_9312_250.n111 a_9312_250.n110 15
R3085 a_9312_250.n144 a_9312_250.n143 15
R3086 a_9312_250.n152 a_9312_250.n151 15
R3087 a_9312_250.n160 a_9312_250.n159 15
R3088 a_9312_250.n168 a_9312_250.n167 15
R3089 a_9312_250.n121 a_9312_250.n120 15
R3090 a_9312_250.n113 a_9312_250.n112 15
R3091 a_9312_250.n141 a_9312_250.n140 15
R3092 a_9312_250.n149 a_9312_250.n148 15
R3093 a_9312_250.n157 a_9312_250.n156 15
R3094 a_9312_250.n165 a_9312_250.n164 15
R3095 a_9312_250.n31 a_9312_250.n30 15
R3096 a_9312_250.n23 a_9312_250.n22 15
R3097 a_9312_250.n15 a_9312_250.n14 15
R3098 a_9312_250.n7 a_9312_250.n6 15
R3099 a_9312_250.n179 a_9312_250.n178 15
R3100 a_9312_250.n39 a_9312_250.n38 15
R3101 a_9312_250.n33 a_9312_250.n32 15
R3102 a_9312_250.n25 a_9312_250.n24 15
R3103 a_9312_250.n17 a_9312_250.n16 15
R3104 a_9312_250.n9 a_9312_250.n8 15
R3105 a_9312_250.n176 a_9312_250.n175 15
R3106 a_9312_250.n122 a_9312_250.n121 14.586
R3107 a_9312_250.n55 a_9312_250.n54 14.523
R3108 a_9312_250.n172 a_9312_250.n171 13.634
R3109 a_9312_250.n183 a_9312_250.n182 13.634
R3110 a_9312_250.n105 a_9312_250.n104 13.624
R3111 a_9312_250.n84 a_9312_250.n83 13.548
R3112 a_9312_250.n47 a_9312_250.n46 12.917
R3113 a_9312_250.n74 a_9312_250.n72 12.917
R3114 a_9312_250.n82 a_9312_250.n80 12.917
R3115 a_9312_250.n90 a_9312_250.n88 12.917
R3116 a_9312_250.n98 a_9312_250.n96 12.917
R3117 a_9312_250.n165 a_9312_250.n163 12.917
R3118 a_9312_250.n157 a_9312_250.n155 12.917
R3119 a_9312_250.n149 a_9312_250.n147 12.917
R3120 a_9312_250.n141 a_9312_250.n139 12.917
R3121 a_9312_250.n114 a_9312_250.n113 12.917
R3122 a_9312_250.n10 a_9312_250.n9 12.917
R3123 a_9312_250.n18 a_9312_250.n17 12.917
R3124 a_9312_250.n26 a_9312_250.n25 12.917
R3125 a_9312_250.n34 a_9312_250.n33 12.917
R3126 a_9312_250.n151 a_9312_250.n150 12.727
R3127 a_9312_250.n14 a_9312_250.n13 12.727
R3128 a_9312_250.n76 a_9312_250.n75 9.677
R3129 a_9312_250.n143 a_9312_250.n142 9.09
R3130 a_9312_250.n22 a_9312_250.n21 9.09
R3131 a_9312_250.n106 a_9312_250.n105 8.708
R3132 a_9312_250.n173 a_9312_250.n172 8.695
R3133 a_9312_250.n184 a_9312_250.n183 8.695
R3134 a_9312_250.n43 a_9312_250.n42 5.806
R3135 a_9312_250.n54 a_9312_250.n52 5.741
R3136 a_9312_250.n48 a_9312_250.n47 5.741
R3137 a_9312_250.n115 a_9312_250.n114 5.741
R3138 a_9312_250.n121 a_9312_250.n119 5.741
R3139 a_9312_250.n35 a_9312_250.n34 5.741
R3140 a_9312_250.n38 a_9312_250.n37 5.741
R3141 a_9312_250.n110 a_9312_250.n109 5.454
R3142 a_9312_250.n30 a_9312_250.n29 5.454
R3143 a_9312_250.n46 a_9312_250.n44 5.023
R3144 a_9312_250.n113 a_9312_250.n111 5.023
R3145 a_9312_250.n27 a_9312_250.n26 5.023
R3146 a_9312_250.n33 a_9312_250.n31 5.023
R3147 a_9312_250.n77 a_9312_250.n74 4.305
R3148 a_9312_250.n80 a_9312_250.n79 4.305
R3149 a_9312_250.n147 a_9312_250.n146 4.305
R3150 a_9312_250.n144 a_9312_250.n141 4.305
R3151 a_9312_250.n19 a_9312_250.n18 4.305
R3152 a_9312_250.n25 a_9312_250.n23 4.305
R3153 a_9312_250.n102 a_9312_250.n101 3.947
R3154 a_9312_250.n103 a_9312_250.n102 3.947
R3155 a_9312_250.n170 a_9312_250.n169 3.947
R3156 a_9312_250.n169 a_9312_250.n168 3.947
R3157 a_9312_250.n181 a_9312_250.n180 3.947
R3158 a_9312_250.n180 a_9312_250.n179 3.947
R3159 a_9312_250.n85 a_9312_250.n82 3.588
R3160 a_9312_250.n88 a_9312_250.n87 3.588
R3161 a_9312_250.n155 a_9312_250.n154 3.588
R3162 a_9312_250.n152 a_9312_250.n149 3.588
R3163 a_9312_250.n11 a_9312_250.n10 3.588
R3164 a_9312_250.n17 a_9312_250.n15 3.588
R3165 a_9312_250.n94 a_9312_250.n93 3.229
R3166 a_9312_250.n95 a_9312_250.n94 3.229
R3167 a_9312_250.n162 a_9312_250.n161 3.229
R3168 a_9312_250.n161 a_9312_250.n160 3.229
R3169 a_9312_250.n4 a_9312_250.n3 3.229
R3170 a_9312_250.n7 a_9312_250.n4 3.229
R3171 a_9312_250.n93 a_9312_250.n90 2.87
R3172 a_9312_250.n96 a_9312_250.n95 2.87
R3173 a_9312_250.n163 a_9312_250.n162 2.87
R3174 a_9312_250.n160 a_9312_250.n157 2.87
R3175 a_9312_250.n3 a_9312_250.n2 2.87
R3176 a_9312_250.n9 a_9312_250.n7 2.87
R3177 a_9312_250.n86 a_9312_250.n85 2.511
R3178 a_9312_250.n87 a_9312_250.n86 2.511
R3179 a_9312_250.n154 a_9312_250.n153 2.511
R3180 a_9312_250.n153 a_9312_250.n152 2.511
R3181 a_9312_250.n12 a_9312_250.n11 2.511
R3182 a_9312_250.n15 a_9312_250.n12 2.511
R3183 a_9312_250.n101 a_9312_250.n98 2.152
R3184 a_9312_250.n104 a_9312_250.n103 2.152
R3185 a_9312_250.n171 a_9312_250.n170 2.152
R3186 a_9312_250.n168 a_9312_250.n165 2.152
R3187 a_9312_250.n182 a_9312_250.n181 2.152
R3188 a_9312_250.n179 a_9312_250.n176 2.152
R3189 a_9312_250.n51 a_9312_250.n50 1.935
R3190 a_9312_250.n118 a_9312_250.n117 1.818
R3191 a_9312_250.n1 a_9312_250.n0 1.818
R3192 a_9312_250.n78 a_9312_250.n77 1.794
R3193 a_9312_250.n79 a_9312_250.n78 1.794
R3194 a_9312_250.n146 a_9312_250.n145 1.794
R3195 a_9312_250.n145 a_9312_250.n144 1.794
R3196 a_9312_250.n20 a_9312_250.n19 1.794
R3197 a_9312_250.n23 a_9312_250.n20 1.794
R3198 a_9312_250.n44 a_9312_250.n41 1.076
R3199 a_9312_250.n41 a_9312_250.n40 1.076
R3200 a_9312_250.n108 a_9312_250.n107 1.076
R3201 a_9312_250.n111 a_9312_250.n108 1.076
R3202 a_9312_250.n28 a_9312_250.n27 1.076
R3203 a_9312_250.n31 a_9312_250.n28 1.076
R3204 a_9312_250.n52 a_9312_250.n49 0.358
R3205 a_9312_250.n49 a_9312_250.n48 0.358
R3206 a_9312_250.n116 a_9312_250.n115 0.358
R3207 a_9312_250.n119 a_9312_250.n116 0.358
R3208 a_9312_250.n36 a_9312_250.n35 0.358
R3209 a_9312_250.n37 a_9312_250.n36 0.358
R3210 a_9312_250.n57 a_9312_250.n56 0.144
R3211 a_9312_250.n60 a_9312_250.n59 0.144
R3212 a_9312_250.n63 a_9312_250.n62 0.144
R3213 a_9312_250.n66 a_9312_250.n65 0.144
R3214 a_9312_250.n69 a_9312_250.n68 0.144
R3215 a_9312_250.n136 a_9312_250.n135 0.144
R3216 a_9312_250.n133 a_9312_250.n132 0.144
R3217 a_9312_250.n130 a_9312_250.n129 0.144
R3218 a_9312_250.n127 a_9312_250.n126 0.144
R3219 a_9312_250.n124 a_9312_250.n123 0.144
R3220 a_9312_250.n59 a_9312_250.n58 0.038
R3221 a_9312_250.n126 a_9312_250.n125 0.038
R3222 a_9312_250.n62 a_9312_250.n61 0.032
R3223 a_9312_250.n129 a_9312_250.n128 0.032
R3224 a_9312_250.n70 a_9312_250.n69 0.029
R3225 a_9312_250.n137 a_9312_250.n136 0.029
R3226 a_9312_250.n65 a_9312_250.n64 0.027
R3227 a_9312_250.n132 a_9312_250.n131 0.027
R3228 a_9312_250.n67 a_9312_250.n66 0.024
R3229 a_9312_250.n134 a_9312_250.n133 0.024
R3230 a_9312_250.n68 a_9312_250.n67 0.021
R3231 a_9312_250.n135 a_9312_250.n134 0.021
R3232 a_9312_250.n64 a_9312_250.n63 0.019
R3233 a_9312_250.n131 a_9312_250.n130 0.019
R3234 a_9312_250.n71 a_9312_250.n70 0.016
R3235 a_9312_250.n138 a_9312_250.n137 0.016
R3236 a_9312_250.n61 a_9312_250.n60 0.013
R3237 a_9312_250.n128 a_9312_250.n127 0.013
R3238 a_9312_250.n58 a_9312_250.n57 0.008
R3239 a_9312_250.n125 a_9312_250.n124 0.008
R3240 a_4490_3828.n45 a_4490_3828.n44 1192.34
R3241 a_4490_3828.n42 a_4490_3828.n41 1031.48
R3242 a_4490_3828.n43 a_4490_3828.t3 1031.48
R3243 a_4490_3828.n117 a_4490_3828.n116 963.661
R3244 a_4490_3828.n119 a_4490_3828.t4 948.736
R3245 a_4490_3828.n42 a_4490_3828.n40 877.239
R3246 a_4490_3828.n44 a_4490_3828.n43 877.239
R3247 a_4490_3828.n118 a_4490_3828.n114 854.746
R3248 a_4490_3828.n117 a_4490_3828.n115 841.893
R3249 a_4490_3828.n120 a_4490_3828.t1 221.779
R3250 a_4490_3828.n45 a_4490_3828.t5 207.807
R3251 a_4490_3828.n113 a_4490_3828.n112 185.223
R3252 a_4490_3828.n120 a_4490_3828.n119 167.141
R3253 a_4490_3828.n131 a_4490_3828.n121 163.552
R3254 a_4490_3828.n43 a_4490_3828.n42 154.24
R3255 a_4490_3828.n118 a_4490_3828.n117 137.116
R3256 a_4490_3828.n61 a_4490_3828.t0 64.755
R3257 a_4490_3828.n112 a_4490_3828.n77 49.503
R3258 a_4490_3828.t2 a_4490_3828.n131 122.225
R3259 a_4490_3828.n106 a_4490_3828.n105 32.833
R3260 a_4490_3828.t2 a_4490_3828.n39 32.727
R3261 a_4490_3828.n62 a_4490_3828.n61 30.598
R3262 a_4490_3828.n39 a_4490_3828.n1 29.09
R3263 a_4490_3828.n98 a_4490_3828.n97 26.863
R3264 a_4490_3828.n119 a_4490_3828.n118 24.1
R3265 a_4490_3828.n90 a_4490_3828.n89 20.893
R3266 a_4490_3828.n125 a_4490_3828.n124 20
R3267 a_4490_3828.n6 a_4490_3828.n5 16.363
R3268 a_4490_3828.n58 a_4490_3828.n57 15
R3269 a_4490_3828.n50 a_4490_3828.n49 15
R3270 a_4490_3828.n83 a_4490_3828.n82 15
R3271 a_4490_3828.n91 a_4490_3828.n90 15
R3272 a_4490_3828.n99 a_4490_3828.n98 15
R3273 a_4490_3828.n60 a_4490_3828.n59 15
R3274 a_4490_3828.n52 a_4490_3828.n51 15
R3275 a_4490_3828.n80 a_4490_3828.n79 15
R3276 a_4490_3828.n88 a_4490_3828.n87 15
R3277 a_4490_3828.n96 a_4490_3828.n95 15
R3278 a_4490_3828.n104 a_4490_3828.n103 15
R3279 a_4490_3828.n107 a_4490_3828.n106 15
R3280 a_4490_3828.n31 a_4490_3828.n30 15
R3281 a_4490_3828.n23 a_4490_3828.n22 15
R3282 a_4490_3828.n15 a_4490_3828.n14 15
R3283 a_4490_3828.n7 a_4490_3828.n6 15
R3284 a_4490_3828.n126 a_4490_3828.n125 15
R3285 a_4490_3828.n39 a_4490_3828.n38 15
R3286 a_4490_3828.n33 a_4490_3828.n32 15
R3287 a_4490_3828.n25 a_4490_3828.n24 15
R3288 a_4490_3828.n17 a_4490_3828.n16 15
R3289 a_4490_3828.n9 a_4490_3828.n8 15
R3290 a_4490_3828.n123 a_4490_3828.n122 15
R3291 a_4490_3828.n82 a_4490_3828.n81 14.924
R3292 a_4490_3828.n61 a_4490_3828.n60 14.123
R3293 a_4490_3828.n130 a_4490_3828.n129 13.634
R3294 a_4490_3828.n111 a_4490_3828.n110 13.544
R3295 a_4490_3828.n53 a_4490_3828.n52 12.917
R3296 a_4490_3828.n80 a_4490_3828.n78 12.917
R3297 a_4490_3828.n88 a_4490_3828.n86 12.917
R3298 a_4490_3828.n96 a_4490_3828.n94 12.917
R3299 a_4490_3828.n104 a_4490_3828.n102 12.917
R3300 a_4490_3828.n10 a_4490_3828.n9 12.917
R3301 a_4490_3828.n18 a_4490_3828.n17 12.917
R3302 a_4490_3828.n26 a_4490_3828.n25 12.917
R3303 a_4490_3828.n34 a_4490_3828.n33 12.917
R3304 a_4490_3828.n14 a_4490_3828.n13 12.727
R3305 a_4490_3828.n113 a_4490_3828.n45 11.069
R3306 a_4490_3828.n22 a_4490_3828.n21 9.09
R3307 a_4490_3828.n49 a_4490_3828.n48 8.954
R3308 a_4490_3828.n112 a_4490_3828.n111 8.805
R3309 a_4490_3828.n131 a_4490_3828.n130 8.695
R3310 a_4490_3828.n60 a_4490_3828.n58 5.741
R3311 a_4490_3828.n54 a_4490_3828.n53 5.741
R3312 a_4490_3828.n35 a_4490_3828.n34 5.741
R3313 a_4490_3828.n38 a_4490_3828.n37 5.741
R3314 a_4490_3828.n30 a_4490_3828.n29 5.454
R3315 a_4490_3828.n52 a_4490_3828.n50 5.023
R3316 a_4490_3828.n27 a_4490_3828.n26 5.023
R3317 a_4490_3828.n33 a_4490_3828.n31 5.023
R3318 a_4490_3828.n83 a_4490_3828.n80 4.305
R3319 a_4490_3828.n86 a_4490_3828.n85 4.305
R3320 a_4490_3828.n19 a_4490_3828.n18 4.305
R3321 a_4490_3828.n25 a_4490_3828.n23 4.305
R3322 a_4490_3828.n108 a_4490_3828.n107 3.947
R3323 a_4490_3828.n109 a_4490_3828.n108 3.947
R3324 a_4490_3828.n128 a_4490_3828.n127 3.947
R3325 a_4490_3828.n127 a_4490_3828.n126 3.947
R3326 a_4490_3828.n91 a_4490_3828.n88 3.588
R3327 a_4490_3828.n94 a_4490_3828.n93 3.588
R3328 a_4490_3828.n11 a_4490_3828.n10 3.588
R3329 a_4490_3828.n17 a_4490_3828.n15 3.588
R3330 a_4490_3828.n100 a_4490_3828.n99 3.229
R3331 a_4490_3828.n101 a_4490_3828.n100 3.229
R3332 a_4490_3828.n4 a_4490_3828.n3 3.229
R3333 a_4490_3828.n7 a_4490_3828.n4 3.229
R3334 a_4490_3828.n57 a_4490_3828.n56 2.984
R3335 a_4490_3828.n99 a_4490_3828.n96 2.87
R3336 a_4490_3828.n102 a_4490_3828.n101 2.87
R3337 a_4490_3828.n3 a_4490_3828.n2 2.87
R3338 a_4490_3828.n9 a_4490_3828.n7 2.87
R3339 a_4490_3828.n92 a_4490_3828.n91 2.511
R3340 a_4490_3828.n93 a_4490_3828.n92 2.511
R3341 a_4490_3828.n12 a_4490_3828.n11 2.511
R3342 a_4490_3828.n15 a_4490_3828.n12 2.511
R3343 a_4490_3828.n107 a_4490_3828.n104 2.152
R3344 a_4490_3828.n110 a_4490_3828.n109 2.152
R3345 a_4490_3828.n129 a_4490_3828.n128 2.152
R3346 a_4490_3828.n126 a_4490_3828.n123 2.152
R3347 a_4490_3828.n1 a_4490_3828.n0 1.818
R3348 a_4490_3828.n84 a_4490_3828.n83 1.794
R3349 a_4490_3828.n85 a_4490_3828.n84 1.794
R3350 a_4490_3828.n20 a_4490_3828.n19 1.794
R3351 a_4490_3828.n23 a_4490_3828.n20 1.794
R3352 a_4490_3828.n121 a_4490_3828.n113 1.165
R3353 a_4490_3828.n50 a_4490_3828.n47 1.076
R3354 a_4490_3828.n47 a_4490_3828.n46 1.076
R3355 a_4490_3828.n28 a_4490_3828.n27 1.076
R3356 a_4490_3828.n31 a_4490_3828.n28 1.076
R3357 a_4490_3828.n121 a_4490_3828.n120 1
R3358 a_4490_3828.n58 a_4490_3828.n55 0.358
R3359 a_4490_3828.n55 a_4490_3828.n54 0.358
R3360 a_4490_3828.n36 a_4490_3828.n35 0.358
R3361 a_4490_3828.n37 a_4490_3828.n36 0.358
R3362 a_4490_3828.n63 a_4490_3828.n62 0.144
R3363 a_4490_3828.n66 a_4490_3828.n65 0.144
R3364 a_4490_3828.n69 a_4490_3828.n68 0.144
R3365 a_4490_3828.n72 a_4490_3828.n71 0.144
R3366 a_4490_3828.n75 a_4490_3828.n74 0.144
R3367 a_4490_3828.n65 a_4490_3828.n64 0.038
R3368 a_4490_3828.n68 a_4490_3828.n67 0.032
R3369 a_4490_3828.n76 a_4490_3828.n75 0.029
R3370 a_4490_3828.n71 a_4490_3828.n70 0.027
R3371 a_4490_3828.n73 a_4490_3828.n72 0.024
R3372 a_4490_3828.n74 a_4490_3828.n73 0.021
R3373 a_4490_3828.n70 a_4490_3828.n69 0.019
R3374 a_4490_3828.n77 a_4490_3828.n76 0.016
R3375 a_4490_3828.n67 a_4490_3828.n66 0.013
R3376 a_4490_3828.n64 a_4490_3828.n63 0.008
R3377 a_3230_5590.n144 a_3230_5590.n143 288.128
R3378 a_3230_5590.n143 a_3230_5590.n142 255.907
R3379 a_3230_5590.n143 a_3230_5590.n75 238.306
R3380 a_3230_5590.n24 a_3230_5590.t0 68.375
R3381 a_3230_5590.n91 a_3230_5590.t2 64.755
R3382 a_3230_5590.t1 a_3230_5590.n199 53.727
R3383 a_3230_5590.n142 a_3230_5590.n107 49.503
R3384 a_3230_5590.n75 a_3230_5590.n40 49.503
R3385 a_3230_5590.n145 a_3230_5590.n144 49.503
R3386 a_3230_5590.n69 a_3230_5590.n68 34.951
R3387 a_3230_5590.n136 a_3230_5590.n135 32.833
R3388 a_3230_5590.n3 a_3230_5590.n2 32.833
R3389 a_3230_5590.n25 a_3230_5590.n24 30.732
R3390 a_3230_5590.n92 a_3230_5590.n91 30.598
R3391 a_3230_5590.t1 a_3230_5590.n159 95.496
R3392 a_3230_5590.n61 a_3230_5590.n60 28.596
R3393 a_3230_5590.n128 a_3230_5590.n127 26.863
R3394 a_3230_5590.n164 a_3230_5590.n163 26.863
R3395 a_3230_5590.n53 a_3230_5590.n52 22.241
R3396 a_3230_5590.n120 a_3230_5590.n119 20.893
R3397 a_3230_5590.n172 a_3230_5590.n171 20.893
R3398 a_3230_5590.n45 a_3230_5590.n44 15.887
R3399 a_3230_5590.n88 a_3230_5590.n87 15
R3400 a_3230_5590.n80 a_3230_5590.n79 15
R3401 a_3230_5590.n113 a_3230_5590.n112 15
R3402 a_3230_5590.n121 a_3230_5590.n120 15
R3403 a_3230_5590.n129 a_3230_5590.n128 15
R3404 a_3230_5590.n90 a_3230_5590.n89 15
R3405 a_3230_5590.n82 a_3230_5590.n81 15
R3406 a_3230_5590.n110 a_3230_5590.n109 15
R3407 a_3230_5590.n118 a_3230_5590.n117 15
R3408 a_3230_5590.n126 a_3230_5590.n125 15
R3409 a_3230_5590.n134 a_3230_5590.n133 15
R3410 a_3230_5590.n137 a_3230_5590.n136 15
R3411 a_3230_5590.n21 a_3230_5590.n20 15
R3412 a_3230_5590.n13 a_3230_5590.n12 15
R3413 a_3230_5590.n46 a_3230_5590.n45 15
R3414 a_3230_5590.n54 a_3230_5590.n53 15
R3415 a_3230_5590.n62 a_3230_5590.n61 15
R3416 a_3230_5590.n70 a_3230_5590.n69 15
R3417 a_3230_5590.n23 a_3230_5590.n22 15
R3418 a_3230_5590.n15 a_3230_5590.n14 15
R3419 a_3230_5590.n43 a_3230_5590.n42 15
R3420 a_3230_5590.n51 a_3230_5590.n50 15
R3421 a_3230_5590.n59 a_3230_5590.n58 15
R3422 a_3230_5590.n67 a_3230_5590.n66 15
R3423 a_3230_5590.n197 a_3230_5590.n196 15
R3424 a_3230_5590.n189 a_3230_5590.n188 15
R3425 a_3230_5590.n181 a_3230_5590.n180 15
R3426 a_3230_5590.n173 a_3230_5590.n172 15
R3427 a_3230_5590.n165 a_3230_5590.n164 15
R3428 a_3230_5590.n199 a_3230_5590.n198 15
R3429 a_3230_5590.n191 a_3230_5590.n190 15
R3430 a_3230_5590.n183 a_3230_5590.n182 15
R3431 a_3230_5590.n175 a_3230_5590.n174 15
R3432 a_3230_5590.n167 a_3230_5590.n166 15
R3433 a_3230_5590.n1 a_3230_5590.n0 15
R3434 a_3230_5590.n4 a_3230_5590.n3 15
R3435 a_3230_5590.n112 a_3230_5590.n111 14.924
R3436 a_3230_5590.n180 a_3230_5590.n179 14.924
R3437 a_3230_5590.n91 a_3230_5590.n90 14.123
R3438 a_3230_5590.n24 a_3230_5590.n23 14.071
R3439 a_3230_5590.n141 a_3230_5590.n140 13.544
R3440 a_3230_5590.n8 a_3230_5590.n7 13.544
R3441 a_3230_5590.n74 a_3230_5590.n73 13.532
R3442 a_3230_5590.n83 a_3230_5590.n82 12.917
R3443 a_3230_5590.n110 a_3230_5590.n108 12.917
R3444 a_3230_5590.n118 a_3230_5590.n116 12.917
R3445 a_3230_5590.n126 a_3230_5590.n124 12.917
R3446 a_3230_5590.n134 a_3230_5590.n132 12.917
R3447 a_3230_5590.n67 a_3230_5590.n65 12.917
R3448 a_3230_5590.n59 a_3230_5590.n57 12.917
R3449 a_3230_5590.n51 a_3230_5590.n49 12.917
R3450 a_3230_5590.n43 a_3230_5590.n41 12.917
R3451 a_3230_5590.n16 a_3230_5590.n15 12.917
R3452 a_3230_5590.n192 a_3230_5590.n191 12.917
R3453 a_3230_5590.n184 a_3230_5590.n183 12.917
R3454 a_3230_5590.n176 a_3230_5590.n175 12.917
R3455 a_3230_5590.n168 a_3230_5590.n167 12.917
R3456 a_3230_5590.n12 a_3230_5590.n11 9.532
R3457 a_3230_5590.n79 a_3230_5590.n78 8.954
R3458 a_3230_5590.n188 a_3230_5590.n187 8.954
R3459 a_3230_5590.n75 a_3230_5590.n74 8.82
R3460 a_3230_5590.n142 a_3230_5590.n141 8.805
R3461 a_3230_5590.n144 a_3230_5590.n8 8.805
R3462 a_3230_5590.n90 a_3230_5590.n88 5.741
R3463 a_3230_5590.n84 a_3230_5590.n83 5.741
R3464 a_3230_5590.n17 a_3230_5590.n16 5.741
R3465 a_3230_5590.n23 a_3230_5590.n21 5.741
R3466 a_3230_5590.n198 a_3230_5590.n197 5.741
R3467 a_3230_5590.n193 a_3230_5590.n192 5.741
R3468 a_3230_5590.n82 a_3230_5590.n80 5.023
R3469 a_3230_5590.n15 a_3230_5590.n13 5.023
R3470 a_3230_5590.n191 a_3230_5590.n189 5.023
R3471 a_3230_5590.n185 a_3230_5590.n184 5.023
R3472 a_3230_5590.n113 a_3230_5590.n110 4.305
R3473 a_3230_5590.n116 a_3230_5590.n115 4.305
R3474 a_3230_5590.n49 a_3230_5590.n48 4.305
R3475 a_3230_5590.n46 a_3230_5590.n43 4.305
R3476 a_3230_5590.n183 a_3230_5590.n181 4.305
R3477 a_3230_5590.n177 a_3230_5590.n176 4.305
R3478 a_3230_5590.n138 a_3230_5590.n137 3.947
R3479 a_3230_5590.n139 a_3230_5590.n138 3.947
R3480 a_3230_5590.n72 a_3230_5590.n71 3.947
R3481 a_3230_5590.n71 a_3230_5590.n70 3.947
R3482 a_3230_5590.n5 a_3230_5590.n4 3.947
R3483 a_3230_5590.n6 a_3230_5590.n5 3.947
R3484 a_3230_5590.n121 a_3230_5590.n118 3.588
R3485 a_3230_5590.n124 a_3230_5590.n123 3.588
R3486 a_3230_5590.n57 a_3230_5590.n56 3.588
R3487 a_3230_5590.n54 a_3230_5590.n51 3.588
R3488 a_3230_5590.n175 a_3230_5590.n173 3.588
R3489 a_3230_5590.n169 a_3230_5590.n168 3.588
R3490 a_3230_5590.n130 a_3230_5590.n129 3.229
R3491 a_3230_5590.n131 a_3230_5590.n130 3.229
R3492 a_3230_5590.n64 a_3230_5590.n63 3.229
R3493 a_3230_5590.n63 a_3230_5590.n62 3.229
R3494 a_3230_5590.n165 a_3230_5590.n162 3.229
R3495 a_3230_5590.n162 a_3230_5590.n161 3.229
R3496 a_3230_5590.n20 a_3230_5590.n19 3.177
R3497 a_3230_5590.n87 a_3230_5590.n86 2.984
R3498 a_3230_5590.n196 a_3230_5590.n195 2.984
R3499 a_3230_5590.n129 a_3230_5590.n126 2.87
R3500 a_3230_5590.n132 a_3230_5590.n131 2.87
R3501 a_3230_5590.n65 a_3230_5590.n64 2.87
R3502 a_3230_5590.n62 a_3230_5590.n59 2.87
R3503 a_3230_5590.n167 a_3230_5590.n165 2.87
R3504 a_3230_5590.n161 a_3230_5590.n160 2.87
R3505 a_3230_5590.n122 a_3230_5590.n121 2.511
R3506 a_3230_5590.n123 a_3230_5590.n122 2.511
R3507 a_3230_5590.n56 a_3230_5590.n55 2.511
R3508 a_3230_5590.n55 a_3230_5590.n54 2.511
R3509 a_3230_5590.n173 a_3230_5590.n170 2.511
R3510 a_3230_5590.n170 a_3230_5590.n169 2.511
R3511 a_3230_5590.n137 a_3230_5590.n134 2.152
R3512 a_3230_5590.n140 a_3230_5590.n139 2.152
R3513 a_3230_5590.n73 a_3230_5590.n72 2.152
R3514 a_3230_5590.n70 a_3230_5590.n67 2.152
R3515 a_3230_5590.n4 a_3230_5590.n1 2.152
R3516 a_3230_5590.n7 a_3230_5590.n6 2.152
R3517 a_3230_5590.n114 a_3230_5590.n113 1.794
R3518 a_3230_5590.n115 a_3230_5590.n114 1.794
R3519 a_3230_5590.n48 a_3230_5590.n47 1.794
R3520 a_3230_5590.n47 a_3230_5590.n46 1.794
R3521 a_3230_5590.n181 a_3230_5590.n178 1.794
R3522 a_3230_5590.n178 a_3230_5590.n177 1.794
R3523 a_3230_5590.n80 a_3230_5590.n77 1.076
R3524 a_3230_5590.n77 a_3230_5590.n76 1.076
R3525 a_3230_5590.n10 a_3230_5590.n9 1.076
R3526 a_3230_5590.n13 a_3230_5590.n10 1.076
R3527 a_3230_5590.n189 a_3230_5590.n186 1.076
R3528 a_3230_5590.n186 a_3230_5590.n185 1.076
R3529 a_3230_5590.n88 a_3230_5590.n85 0.358
R3530 a_3230_5590.n85 a_3230_5590.n84 0.358
R3531 a_3230_5590.n18 a_3230_5590.n17 0.358
R3532 a_3230_5590.n21 a_3230_5590.n18 0.358
R3533 a_3230_5590.n197 a_3230_5590.n194 0.358
R3534 a_3230_5590.n194 a_3230_5590.n193 0.358
R3535 a_3230_5590.n93 a_3230_5590.n92 0.144
R3536 a_3230_5590.n96 a_3230_5590.n95 0.144
R3537 a_3230_5590.n99 a_3230_5590.n98 0.144
R3538 a_3230_5590.n102 a_3230_5590.n101 0.144
R3539 a_3230_5590.n105 a_3230_5590.n104 0.144
R3540 a_3230_5590.n38 a_3230_5590.n37 0.144
R3541 a_3230_5590.n35 a_3230_5590.n34 0.144
R3542 a_3230_5590.n32 a_3230_5590.n31 0.144
R3543 a_3230_5590.n29 a_3230_5590.n28 0.144
R3544 a_3230_5590.n26 a_3230_5590.n25 0.144
R3545 a_3230_5590.n157 a_3230_5590.n156 0.144
R3546 a_3230_5590.n154 a_3230_5590.n153 0.144
R3547 a_3230_5590.n151 a_3230_5590.n150 0.144
R3548 a_3230_5590.n148 a_3230_5590.n147 0.144
R3549 a_3230_5590.n95 a_3230_5590.n94 0.038
R3550 a_3230_5590.n28 a_3230_5590.n27 0.038
R3551 a_3230_5590.n158 a_3230_5590.n157 0.038
R3552 a_3230_5590.n98 a_3230_5590.n97 0.032
R3553 a_3230_5590.n31 a_3230_5590.n30 0.032
R3554 a_3230_5590.n155 a_3230_5590.n154 0.032
R3555 a_3230_5590.n106 a_3230_5590.n105 0.029
R3556 a_3230_5590.n39 a_3230_5590.n38 0.029
R3557 a_3230_5590.n147 a_3230_5590.n146 0.029
R3558 a_3230_5590.n101 a_3230_5590.n100 0.027
R3559 a_3230_5590.n34 a_3230_5590.n33 0.027
R3560 a_3230_5590.n152 a_3230_5590.n151 0.027
R3561 a_3230_5590.n103 a_3230_5590.n102 0.024
R3562 a_3230_5590.n36 a_3230_5590.n35 0.024
R3563 a_3230_5590.n150 a_3230_5590.n149 0.024
R3564 a_3230_5590.n104 a_3230_5590.n103 0.021
R3565 a_3230_5590.n37 a_3230_5590.n36 0.021
R3566 a_3230_5590.n149 a_3230_5590.n148 0.021
R3567 a_3230_5590.n100 a_3230_5590.n99 0.019
R3568 a_3230_5590.n33 a_3230_5590.n32 0.019
R3569 a_3230_5590.n153 a_3230_5590.n152 0.019
R3570 a_3230_5590.n107 a_3230_5590.n106 0.016
R3571 a_3230_5590.n40 a_3230_5590.n39 0.016
R3572 a_3230_5590.n146 a_3230_5590.n145 0.016
R3573 a_3230_5590.n97 a_3230_5590.n96 0.013
R3574 a_3230_5590.n30 a_3230_5590.n29 0.013
R3575 a_3230_5590.n156 a_3230_5590.n155 0.013
R3576 a_3230_5590.n94 a_3230_5590.n93 0.008
R3577 a_3230_5590.n27 a_3230_5590.n26 0.008
R3578 a_3230_5590.n159 a_3230_5590.n158 0.008
R3579 a_n1698_2236.n115 a_n1698_2236.n114 1119.08
R3580 a_n1698_2236.n118 a_n1698_2236.n30 1116.79
R3581 a_n1698_2236.n116 a_n1698_2236.n72 1116.76
R3582 a_n1698_2236.n117 a_n1698_2236.n51 1116.76
R3583 a_n1698_2236.n115 a_n1698_2236.n93 1116.75
R3584 a_n1698_2236.n104 a_n1698_2236.t5 1018.63
R3585 a_n1698_2236.n114 a_n1698_2236.n113 1018.63
R3586 a_n1698_2236.n83 a_n1698_2236.n82 1018.63
R3587 a_n1698_2236.n93 a_n1698_2236.n92 1018.63
R3588 a_n1698_2236.n62 a_n1698_2236.t3 1018.63
R3589 a_n1698_2236.n72 a_n1698_2236.n71 1018.63
R3590 a_n1698_2236.n41 a_n1698_2236.t6 1018.63
R3591 a_n1698_2236.n51 a_n1698_2236.n50 1018.63
R3592 a_n1698_2236.n20 a_n1698_2236.n19 1018.63
R3593 a_n1698_2236.n30 a_n1698_2236.n29 1018.63
R3594 a_n1698_2236.n113 a_n1698_2236.n94 864.386
R3595 a_n1698_2236.n112 a_n1698_2236.n95 864.386
R3596 a_n1698_2236.n111 a_n1698_2236.n96 864.386
R3597 a_n1698_2236.n110 a_n1698_2236.n97 864.386
R3598 a_n1698_2236.n109 a_n1698_2236.n98 864.386
R3599 a_n1698_2236.n108 a_n1698_2236.n99 864.386
R3600 a_n1698_2236.n107 a_n1698_2236.n100 864.386
R3601 a_n1698_2236.n106 a_n1698_2236.n101 864.386
R3602 a_n1698_2236.n105 a_n1698_2236.n102 864.386
R3603 a_n1698_2236.n104 a_n1698_2236.n103 864.386
R3604 a_n1698_2236.n92 a_n1698_2236.n73 864.386
R3605 a_n1698_2236.n91 a_n1698_2236.n74 864.386
R3606 a_n1698_2236.n90 a_n1698_2236.n75 864.386
R3607 a_n1698_2236.n89 a_n1698_2236.n76 864.386
R3608 a_n1698_2236.n88 a_n1698_2236.n77 864.386
R3609 a_n1698_2236.n87 a_n1698_2236.n78 864.386
R3610 a_n1698_2236.n86 a_n1698_2236.n79 864.386
R3611 a_n1698_2236.n85 a_n1698_2236.t4 864.386
R3612 a_n1698_2236.n84 a_n1698_2236.n80 864.386
R3613 a_n1698_2236.n83 a_n1698_2236.n81 864.386
R3614 a_n1698_2236.n71 a_n1698_2236.n52 864.386
R3615 a_n1698_2236.n70 a_n1698_2236.n53 864.386
R3616 a_n1698_2236.n69 a_n1698_2236.n54 864.386
R3617 a_n1698_2236.n68 a_n1698_2236.n55 864.386
R3618 a_n1698_2236.n67 a_n1698_2236.n56 864.386
R3619 a_n1698_2236.n66 a_n1698_2236.n57 864.386
R3620 a_n1698_2236.n65 a_n1698_2236.n58 864.386
R3621 a_n1698_2236.n64 a_n1698_2236.n59 864.386
R3622 a_n1698_2236.n63 a_n1698_2236.n60 864.386
R3623 a_n1698_2236.n62 a_n1698_2236.n61 864.386
R3624 a_n1698_2236.n50 a_n1698_2236.n31 864.386
R3625 a_n1698_2236.n49 a_n1698_2236.n32 864.386
R3626 a_n1698_2236.n48 a_n1698_2236.n33 864.386
R3627 a_n1698_2236.n47 a_n1698_2236.n34 864.386
R3628 a_n1698_2236.n46 a_n1698_2236.n35 864.386
R3629 a_n1698_2236.n45 a_n1698_2236.n36 864.386
R3630 a_n1698_2236.n44 a_n1698_2236.n37 864.386
R3631 a_n1698_2236.n43 a_n1698_2236.n38 864.386
R3632 a_n1698_2236.n42 a_n1698_2236.n39 864.386
R3633 a_n1698_2236.n41 a_n1698_2236.n40 864.386
R3634 a_n1698_2236.n29 a_n1698_2236.n10 864.386
R3635 a_n1698_2236.n28 a_n1698_2236.n11 864.386
R3636 a_n1698_2236.n27 a_n1698_2236.n12 864.386
R3637 a_n1698_2236.n26 a_n1698_2236.t7 864.386
R3638 a_n1698_2236.n25 a_n1698_2236.n13 864.386
R3639 a_n1698_2236.n24 a_n1698_2236.n14 864.386
R3640 a_n1698_2236.n23 a_n1698_2236.n15 864.386
R3641 a_n1698_2236.n22 a_n1698_2236.n16 864.386
R3642 a_n1698_2236.n21 a_n1698_2236.n17 864.386
R3643 a_n1698_2236.n20 a_n1698_2236.n18 864.386
R3644 a_n1698_2236.n127 a_n1698_2236.n126 809.76
R3645 a_n1698_2236.n127 a_n1698_2236.n125 691.67
R3646 a_n1698_2236.n128 a_n1698_2236.n124 691.67
R3647 a_n1698_2236.n129 a_n1698_2236.n123 691.67
R3648 a_n1698_2236.n130 a_n1698_2236.n122 691.67
R3649 a_n1698_2236.n131 a_n1698_2236.n121 691.67
R3650 a_n1698_2236.n120 a_n1698_2236.t0 691.67
R3651 a_n1698_2236.n119 a_n1698_2236.n9 691.67
R3652 a_n1698_2236.n148 a_n1698_2236.n147 331.687
R3653 a_n1698_2236.n119 a_n1698_2236.n118 258.096
R3654 a_n1698_2236.n105 a_n1698_2236.n104 154.24
R3655 a_n1698_2236.n106 a_n1698_2236.n105 154.24
R3656 a_n1698_2236.n107 a_n1698_2236.n106 154.24
R3657 a_n1698_2236.n108 a_n1698_2236.n107 154.24
R3658 a_n1698_2236.n109 a_n1698_2236.n108 154.24
R3659 a_n1698_2236.n110 a_n1698_2236.n109 154.24
R3660 a_n1698_2236.n111 a_n1698_2236.n110 154.24
R3661 a_n1698_2236.n112 a_n1698_2236.n111 154.24
R3662 a_n1698_2236.n113 a_n1698_2236.n112 154.24
R3663 a_n1698_2236.n84 a_n1698_2236.n83 154.24
R3664 a_n1698_2236.n85 a_n1698_2236.n84 154.24
R3665 a_n1698_2236.n86 a_n1698_2236.n85 154.24
R3666 a_n1698_2236.n87 a_n1698_2236.n86 154.24
R3667 a_n1698_2236.n88 a_n1698_2236.n87 154.24
R3668 a_n1698_2236.n89 a_n1698_2236.n88 154.24
R3669 a_n1698_2236.n90 a_n1698_2236.n89 154.24
R3670 a_n1698_2236.n91 a_n1698_2236.n90 154.24
R3671 a_n1698_2236.n92 a_n1698_2236.n91 154.24
R3672 a_n1698_2236.n63 a_n1698_2236.n62 154.24
R3673 a_n1698_2236.n64 a_n1698_2236.n63 154.24
R3674 a_n1698_2236.n65 a_n1698_2236.n64 154.24
R3675 a_n1698_2236.n66 a_n1698_2236.n65 154.24
R3676 a_n1698_2236.n67 a_n1698_2236.n66 154.24
R3677 a_n1698_2236.n68 a_n1698_2236.n67 154.24
R3678 a_n1698_2236.n69 a_n1698_2236.n68 154.24
R3679 a_n1698_2236.n70 a_n1698_2236.n69 154.24
R3680 a_n1698_2236.n71 a_n1698_2236.n70 154.24
R3681 a_n1698_2236.n42 a_n1698_2236.n41 154.24
R3682 a_n1698_2236.n43 a_n1698_2236.n42 154.24
R3683 a_n1698_2236.n44 a_n1698_2236.n43 154.24
R3684 a_n1698_2236.n45 a_n1698_2236.n44 154.24
R3685 a_n1698_2236.n46 a_n1698_2236.n45 154.24
R3686 a_n1698_2236.n47 a_n1698_2236.n46 154.24
R3687 a_n1698_2236.n48 a_n1698_2236.n47 154.24
R3688 a_n1698_2236.n49 a_n1698_2236.n48 154.24
R3689 a_n1698_2236.n50 a_n1698_2236.n49 154.24
R3690 a_n1698_2236.n21 a_n1698_2236.n20 154.24
R3691 a_n1698_2236.n22 a_n1698_2236.n21 154.24
R3692 a_n1698_2236.n23 a_n1698_2236.n22 154.24
R3693 a_n1698_2236.n24 a_n1698_2236.n23 154.24
R3694 a_n1698_2236.n25 a_n1698_2236.n24 154.24
R3695 a_n1698_2236.n26 a_n1698_2236.n25 154.24
R3696 a_n1698_2236.n27 a_n1698_2236.n26 154.24
R3697 a_n1698_2236.n28 a_n1698_2236.n27 154.24
R3698 a_n1698_2236.n29 a_n1698_2236.n28 154.24
R3699 a_n1698_2236.n145 a_n1698_2236.n144 121.919
R3700 a_n1698_2236.n138 a_n1698_2236.n137 121.919
R3701 a_n1698_2236.n147 a_n1698_2236.n132 119.693
R3702 a_n1698_2236.n120 a_n1698_2236.n119 118.09
R3703 a_n1698_2236.n131 a_n1698_2236.n130 118.09
R3704 a_n1698_2236.n130 a_n1698_2236.n129 118.09
R3705 a_n1698_2236.n129 a_n1698_2236.n128 118.09
R3706 a_n1698_2236.n128 a_n1698_2236.n127 118.09
R3707 a_n1698_2236.n146 a_n1698_2236.n145 68.894
R3708 a_n1698_2236.n147 a_n1698_2236.n146 68.534
R3709 a_n1698_2236.n132 a_n1698_2236.n131 60.25
R3710 a_n1698_2236.n132 a_n1698_2236.n120 57.84
R3711 a_n1698_2236.n145 a_n1698_2236.n141 51.59
R3712 a_n1698_2236.n138 a_n1698_2236.n135 51.59
R3713 a_n1698_2236.n149 a_n1698_2236.n148 49.503
R3714 a_n1698_2236.t2 a_n1698_2236.n203 32.727
R3715 a_n1698_2236.t2 a_n1698_2236.n163 71.919
R3716 a_n1698_2236.n203 a_n1698_2236.n165 29.09
R3717 a_n1698_2236.n3 a_n1698_2236.n2 20
R3718 a_n1698_2236.n170 a_n1698_2236.n169 16.363
R3719 a_n1698_2236.n195 a_n1698_2236.n194 15
R3720 a_n1698_2236.n187 a_n1698_2236.n186 15
R3721 a_n1698_2236.n179 a_n1698_2236.n178 15
R3722 a_n1698_2236.n171 a_n1698_2236.n170 15
R3723 a_n1698_2236.n203 a_n1698_2236.n202 15
R3724 a_n1698_2236.n197 a_n1698_2236.n196 15
R3725 a_n1698_2236.n189 a_n1698_2236.n188 15
R3726 a_n1698_2236.n181 a_n1698_2236.n180 15
R3727 a_n1698_2236.n173 a_n1698_2236.n172 15
R3728 a_n1698_2236.n1 a_n1698_2236.n0 15
R3729 a_n1698_2236.n4 a_n1698_2236.n3 15
R3730 a_n1698_2236.n8 a_n1698_2236.n7 13.634
R3731 a_n1698_2236.n198 a_n1698_2236.n197 12.917
R3732 a_n1698_2236.n190 a_n1698_2236.n189 12.917
R3733 a_n1698_2236.n182 a_n1698_2236.n181 12.917
R3734 a_n1698_2236.n174 a_n1698_2236.n173 12.917
R3735 a_n1698_2236.n178 a_n1698_2236.n177 12.727
R3736 a_n1698_2236.n186 a_n1698_2236.n185 9.09
R3737 a_n1698_2236.n148 a_n1698_2236.n8 8.695
R3738 a_n1698_2236.n202 a_n1698_2236.n201 5.741
R3739 a_n1698_2236.n199 a_n1698_2236.n198 5.741
R3740 a_n1698_2236.n194 a_n1698_2236.n193 5.454
R3741 a_n1698_2236.n197 a_n1698_2236.n195 5.023
R3742 a_n1698_2236.n191 a_n1698_2236.n190 5.023
R3743 a_n1698_2236.n189 a_n1698_2236.n187 4.305
R3744 a_n1698_2236.n183 a_n1698_2236.n182 4.305
R3745 a_n1698_2236.n5 a_n1698_2236.n4 3.947
R3746 a_n1698_2236.n6 a_n1698_2236.n5 3.947
R3747 a_n1698_2236.n181 a_n1698_2236.n179 3.588
R3748 a_n1698_2236.n175 a_n1698_2236.n174 3.588
R3749 a_n1698_2236.n144 a_n1698_2236.n142 3.48
R3750 a_n1698_2236.n144 a_n1698_2236.n143 3.48
R3751 a_n1698_2236.n141 a_n1698_2236.n139 3.48
R3752 a_n1698_2236.n141 a_n1698_2236.n140 3.48
R3753 a_n1698_2236.n135 a_n1698_2236.n133 3.48
R3754 a_n1698_2236.n135 a_n1698_2236.n134 3.48
R3755 a_n1698_2236.n137 a_n1698_2236.n136 3.48
R3756 a_n1698_2236.n137 a_n1698_2236.t1 3.48
R3757 a_n1698_2236.n171 a_n1698_2236.n168 3.229
R3758 a_n1698_2236.n168 a_n1698_2236.n167 3.229
R3759 a_n1698_2236.n173 a_n1698_2236.n171 2.87
R3760 a_n1698_2236.n167 a_n1698_2236.n166 2.87
R3761 a_n1698_2236.n179 a_n1698_2236.n176 2.511
R3762 a_n1698_2236.n176 a_n1698_2236.n175 2.511
R3763 a_n1698_2236.n116 a_n1698_2236.n115 2.506
R3764 a_n1698_2236.n117 a_n1698_2236.n116 2.457
R3765 a_n1698_2236.n118 a_n1698_2236.n117 2.399
R3766 a_n1698_2236.n4 a_n1698_2236.n1 2.152
R3767 a_n1698_2236.n7 a_n1698_2236.n6 2.152
R3768 a_n1698_2236.n165 a_n1698_2236.n164 1.818
R3769 a_n1698_2236.n187 a_n1698_2236.n184 1.794
R3770 a_n1698_2236.n184 a_n1698_2236.n183 1.794
R3771 a_n1698_2236.n146 a_n1698_2236.n138 1.435
R3772 a_n1698_2236.n195 a_n1698_2236.n192 1.076
R3773 a_n1698_2236.n192 a_n1698_2236.n191 1.076
R3774 a_n1698_2236.n201 a_n1698_2236.n200 0.358
R3775 a_n1698_2236.n200 a_n1698_2236.n199 0.358
R3776 a_n1698_2236.n161 a_n1698_2236.n160 0.144
R3777 a_n1698_2236.n158 a_n1698_2236.n157 0.144
R3778 a_n1698_2236.n155 a_n1698_2236.n154 0.144
R3779 a_n1698_2236.n152 a_n1698_2236.n151 0.144
R3780 a_n1698_2236.n162 a_n1698_2236.n161 0.038
R3781 a_n1698_2236.n159 a_n1698_2236.n158 0.032
R3782 a_n1698_2236.n151 a_n1698_2236.n150 0.029
R3783 a_n1698_2236.n156 a_n1698_2236.n155 0.027
R3784 a_n1698_2236.n154 a_n1698_2236.n153 0.024
R3785 a_n1698_2236.n153 a_n1698_2236.n152 0.021
R3786 a_n1698_2236.n157 a_n1698_2236.n156 0.019
R3787 a_n1698_2236.n150 a_n1698_2236.n149 0.016
R3788 a_n1698_2236.n160 a_n1698_2236.n159 0.013
R3789 a_n1698_2236.n163 a_n1698_2236.n162 0.008
R3790 a_12504_5562.n144 a_12504_5562.n143 297.845
R3791 a_12504_5562.n143 a_12504_5562.n142 255.585
R3792 a_12504_5562.n143 a_12504_5562.n75 169.38
R3793 a_12504_5562.n91 a_12504_5562.t1 64.755
R3794 a_12504_5562.n24 a_12504_5562.t2 64.755
R3795 a_12504_5562.t0 a_12504_5562.n199 53.727
R3796 a_12504_5562.n142 a_12504_5562.n107 49.503
R3797 a_12504_5562.n75 a_12504_5562.n40 49.503
R3798 a_12504_5562.n145 a_12504_5562.n144 49.503
R3799 a_12504_5562.n136 a_12504_5562.n135 32.833
R3800 a_12504_5562.n69 a_12504_5562.n68 32.833
R3801 a_12504_5562.n3 a_12504_5562.n2 32.833
R3802 a_12504_5562.n25 a_12504_5562.n24 30.598
R3803 a_12504_5562.n92 a_12504_5562.n91 30.598
R3804 a_12504_5562.t0 a_12504_5562.n159 95.496
R3805 a_12504_5562.n128 a_12504_5562.n127 26.863
R3806 a_12504_5562.n61 a_12504_5562.n60 26.863
R3807 a_12504_5562.n164 a_12504_5562.n163 26.863
R3808 a_12504_5562.n120 a_12504_5562.n119 20.893
R3809 a_12504_5562.n53 a_12504_5562.n52 20.893
R3810 a_12504_5562.n172 a_12504_5562.n171 20.893
R3811 a_12504_5562.n88 a_12504_5562.n87 15
R3812 a_12504_5562.n80 a_12504_5562.n79 15
R3813 a_12504_5562.n113 a_12504_5562.n112 15
R3814 a_12504_5562.n121 a_12504_5562.n120 15
R3815 a_12504_5562.n129 a_12504_5562.n128 15
R3816 a_12504_5562.n90 a_12504_5562.n89 15
R3817 a_12504_5562.n82 a_12504_5562.n81 15
R3818 a_12504_5562.n110 a_12504_5562.n109 15
R3819 a_12504_5562.n118 a_12504_5562.n117 15
R3820 a_12504_5562.n126 a_12504_5562.n125 15
R3821 a_12504_5562.n134 a_12504_5562.n133 15
R3822 a_12504_5562.n137 a_12504_5562.n136 15
R3823 a_12504_5562.n21 a_12504_5562.n20 15
R3824 a_12504_5562.n13 a_12504_5562.n12 15
R3825 a_12504_5562.n46 a_12504_5562.n45 15
R3826 a_12504_5562.n54 a_12504_5562.n53 15
R3827 a_12504_5562.n62 a_12504_5562.n61 15
R3828 a_12504_5562.n70 a_12504_5562.n69 15
R3829 a_12504_5562.n23 a_12504_5562.n22 15
R3830 a_12504_5562.n15 a_12504_5562.n14 15
R3831 a_12504_5562.n43 a_12504_5562.n42 15
R3832 a_12504_5562.n51 a_12504_5562.n50 15
R3833 a_12504_5562.n59 a_12504_5562.n58 15
R3834 a_12504_5562.n67 a_12504_5562.n66 15
R3835 a_12504_5562.n197 a_12504_5562.n196 15
R3836 a_12504_5562.n189 a_12504_5562.n188 15
R3837 a_12504_5562.n181 a_12504_5562.n180 15
R3838 a_12504_5562.n173 a_12504_5562.n172 15
R3839 a_12504_5562.n165 a_12504_5562.n164 15
R3840 a_12504_5562.n199 a_12504_5562.n198 15
R3841 a_12504_5562.n191 a_12504_5562.n190 15
R3842 a_12504_5562.n183 a_12504_5562.n182 15
R3843 a_12504_5562.n175 a_12504_5562.n174 15
R3844 a_12504_5562.n167 a_12504_5562.n166 15
R3845 a_12504_5562.n1 a_12504_5562.n0 15
R3846 a_12504_5562.n4 a_12504_5562.n3 15
R3847 a_12504_5562.n112 a_12504_5562.n111 14.924
R3848 a_12504_5562.n45 a_12504_5562.n44 14.924
R3849 a_12504_5562.n180 a_12504_5562.n179 14.924
R3850 a_12504_5562.n91 a_12504_5562.n90 14.123
R3851 a_12504_5562.n24 a_12504_5562.n23 14.123
R3852 a_12504_5562.n141 a_12504_5562.n140 13.544
R3853 a_12504_5562.n74 a_12504_5562.n73 13.544
R3854 a_12504_5562.n8 a_12504_5562.n7 13.544
R3855 a_12504_5562.n83 a_12504_5562.n82 12.917
R3856 a_12504_5562.n110 a_12504_5562.n108 12.917
R3857 a_12504_5562.n118 a_12504_5562.n116 12.917
R3858 a_12504_5562.n126 a_12504_5562.n124 12.917
R3859 a_12504_5562.n134 a_12504_5562.n132 12.917
R3860 a_12504_5562.n67 a_12504_5562.n65 12.917
R3861 a_12504_5562.n59 a_12504_5562.n57 12.917
R3862 a_12504_5562.n51 a_12504_5562.n49 12.917
R3863 a_12504_5562.n43 a_12504_5562.n41 12.917
R3864 a_12504_5562.n16 a_12504_5562.n15 12.917
R3865 a_12504_5562.n192 a_12504_5562.n191 12.917
R3866 a_12504_5562.n184 a_12504_5562.n183 12.917
R3867 a_12504_5562.n176 a_12504_5562.n175 12.917
R3868 a_12504_5562.n168 a_12504_5562.n167 12.917
R3869 a_12504_5562.n79 a_12504_5562.n78 8.954
R3870 a_12504_5562.n12 a_12504_5562.n11 8.954
R3871 a_12504_5562.n188 a_12504_5562.n187 8.954
R3872 a_12504_5562.n142 a_12504_5562.n141 8.805
R3873 a_12504_5562.n75 a_12504_5562.n74 8.805
R3874 a_12504_5562.n144 a_12504_5562.n8 8.805
R3875 a_12504_5562.n90 a_12504_5562.n88 5.741
R3876 a_12504_5562.n84 a_12504_5562.n83 5.741
R3877 a_12504_5562.n17 a_12504_5562.n16 5.741
R3878 a_12504_5562.n23 a_12504_5562.n21 5.741
R3879 a_12504_5562.n198 a_12504_5562.n197 5.741
R3880 a_12504_5562.n193 a_12504_5562.n192 5.741
R3881 a_12504_5562.n82 a_12504_5562.n80 5.023
R3882 a_12504_5562.n15 a_12504_5562.n13 5.023
R3883 a_12504_5562.n191 a_12504_5562.n189 5.023
R3884 a_12504_5562.n185 a_12504_5562.n184 5.023
R3885 a_12504_5562.n113 a_12504_5562.n110 4.305
R3886 a_12504_5562.n116 a_12504_5562.n115 4.305
R3887 a_12504_5562.n49 a_12504_5562.n48 4.305
R3888 a_12504_5562.n46 a_12504_5562.n43 4.305
R3889 a_12504_5562.n183 a_12504_5562.n181 4.305
R3890 a_12504_5562.n177 a_12504_5562.n176 4.305
R3891 a_12504_5562.n138 a_12504_5562.n137 3.947
R3892 a_12504_5562.n139 a_12504_5562.n138 3.947
R3893 a_12504_5562.n72 a_12504_5562.n71 3.947
R3894 a_12504_5562.n71 a_12504_5562.n70 3.947
R3895 a_12504_5562.n5 a_12504_5562.n4 3.947
R3896 a_12504_5562.n6 a_12504_5562.n5 3.947
R3897 a_12504_5562.n121 a_12504_5562.n118 3.588
R3898 a_12504_5562.n124 a_12504_5562.n123 3.588
R3899 a_12504_5562.n57 a_12504_5562.n56 3.588
R3900 a_12504_5562.n54 a_12504_5562.n51 3.588
R3901 a_12504_5562.n175 a_12504_5562.n173 3.588
R3902 a_12504_5562.n169 a_12504_5562.n168 3.588
R3903 a_12504_5562.n130 a_12504_5562.n129 3.229
R3904 a_12504_5562.n131 a_12504_5562.n130 3.229
R3905 a_12504_5562.n64 a_12504_5562.n63 3.229
R3906 a_12504_5562.n63 a_12504_5562.n62 3.229
R3907 a_12504_5562.n165 a_12504_5562.n162 3.229
R3908 a_12504_5562.n162 a_12504_5562.n161 3.229
R3909 a_12504_5562.n87 a_12504_5562.n86 2.984
R3910 a_12504_5562.n20 a_12504_5562.n19 2.984
R3911 a_12504_5562.n196 a_12504_5562.n195 2.984
R3912 a_12504_5562.n129 a_12504_5562.n126 2.87
R3913 a_12504_5562.n132 a_12504_5562.n131 2.87
R3914 a_12504_5562.n65 a_12504_5562.n64 2.87
R3915 a_12504_5562.n62 a_12504_5562.n59 2.87
R3916 a_12504_5562.n167 a_12504_5562.n165 2.87
R3917 a_12504_5562.n161 a_12504_5562.n160 2.87
R3918 a_12504_5562.n122 a_12504_5562.n121 2.511
R3919 a_12504_5562.n123 a_12504_5562.n122 2.511
R3920 a_12504_5562.n56 a_12504_5562.n55 2.511
R3921 a_12504_5562.n55 a_12504_5562.n54 2.511
R3922 a_12504_5562.n173 a_12504_5562.n170 2.511
R3923 a_12504_5562.n170 a_12504_5562.n169 2.511
R3924 a_12504_5562.n137 a_12504_5562.n134 2.152
R3925 a_12504_5562.n140 a_12504_5562.n139 2.152
R3926 a_12504_5562.n73 a_12504_5562.n72 2.152
R3927 a_12504_5562.n70 a_12504_5562.n67 2.152
R3928 a_12504_5562.n4 a_12504_5562.n1 2.152
R3929 a_12504_5562.n7 a_12504_5562.n6 2.152
R3930 a_12504_5562.n114 a_12504_5562.n113 1.794
R3931 a_12504_5562.n115 a_12504_5562.n114 1.794
R3932 a_12504_5562.n48 a_12504_5562.n47 1.794
R3933 a_12504_5562.n47 a_12504_5562.n46 1.794
R3934 a_12504_5562.n181 a_12504_5562.n178 1.794
R3935 a_12504_5562.n178 a_12504_5562.n177 1.794
R3936 a_12504_5562.n80 a_12504_5562.n77 1.076
R3937 a_12504_5562.n77 a_12504_5562.n76 1.076
R3938 a_12504_5562.n10 a_12504_5562.n9 1.076
R3939 a_12504_5562.n13 a_12504_5562.n10 1.076
R3940 a_12504_5562.n189 a_12504_5562.n186 1.076
R3941 a_12504_5562.n186 a_12504_5562.n185 1.076
R3942 a_12504_5562.n88 a_12504_5562.n85 0.358
R3943 a_12504_5562.n85 a_12504_5562.n84 0.358
R3944 a_12504_5562.n18 a_12504_5562.n17 0.358
R3945 a_12504_5562.n21 a_12504_5562.n18 0.358
R3946 a_12504_5562.n197 a_12504_5562.n194 0.358
R3947 a_12504_5562.n194 a_12504_5562.n193 0.358
R3948 a_12504_5562.n93 a_12504_5562.n92 0.144
R3949 a_12504_5562.n96 a_12504_5562.n95 0.144
R3950 a_12504_5562.n99 a_12504_5562.n98 0.144
R3951 a_12504_5562.n102 a_12504_5562.n101 0.144
R3952 a_12504_5562.n105 a_12504_5562.n104 0.144
R3953 a_12504_5562.n38 a_12504_5562.n37 0.144
R3954 a_12504_5562.n35 a_12504_5562.n34 0.144
R3955 a_12504_5562.n32 a_12504_5562.n31 0.144
R3956 a_12504_5562.n29 a_12504_5562.n28 0.144
R3957 a_12504_5562.n26 a_12504_5562.n25 0.144
R3958 a_12504_5562.n157 a_12504_5562.n156 0.144
R3959 a_12504_5562.n154 a_12504_5562.n153 0.144
R3960 a_12504_5562.n151 a_12504_5562.n150 0.144
R3961 a_12504_5562.n148 a_12504_5562.n147 0.144
R3962 a_12504_5562.n95 a_12504_5562.n94 0.038
R3963 a_12504_5562.n28 a_12504_5562.n27 0.038
R3964 a_12504_5562.n158 a_12504_5562.n157 0.038
R3965 a_12504_5562.n98 a_12504_5562.n97 0.032
R3966 a_12504_5562.n31 a_12504_5562.n30 0.032
R3967 a_12504_5562.n155 a_12504_5562.n154 0.032
R3968 a_12504_5562.n106 a_12504_5562.n105 0.029
R3969 a_12504_5562.n39 a_12504_5562.n38 0.029
R3970 a_12504_5562.n147 a_12504_5562.n146 0.029
R3971 a_12504_5562.n101 a_12504_5562.n100 0.027
R3972 a_12504_5562.n34 a_12504_5562.n33 0.027
R3973 a_12504_5562.n152 a_12504_5562.n151 0.027
R3974 a_12504_5562.n103 a_12504_5562.n102 0.024
R3975 a_12504_5562.n36 a_12504_5562.n35 0.024
R3976 a_12504_5562.n150 a_12504_5562.n149 0.024
R3977 a_12504_5562.n104 a_12504_5562.n103 0.021
R3978 a_12504_5562.n37 a_12504_5562.n36 0.021
R3979 a_12504_5562.n149 a_12504_5562.n148 0.021
R3980 a_12504_5562.n100 a_12504_5562.n99 0.019
R3981 a_12504_5562.n33 a_12504_5562.n32 0.019
R3982 a_12504_5562.n153 a_12504_5562.n152 0.019
R3983 a_12504_5562.n107 a_12504_5562.n106 0.016
R3984 a_12504_5562.n40 a_12504_5562.n39 0.016
R3985 a_12504_5562.n146 a_12504_5562.n145 0.016
R3986 a_12504_5562.n97 a_12504_5562.n96 0.013
R3987 a_12504_5562.n30 a_12504_5562.n29 0.013
R3988 a_12504_5562.n156 a_12504_5562.n155 0.013
R3989 a_12504_5562.n94 a_12504_5562.n93 0.008
R3990 a_12504_5562.n27 a_12504_5562.n26 0.008
R3991 a_12504_5562.n159 a_12504_5562.n158 0.008
R3992 OUT.n147 OUT.n146 1369.18
R3993 OUT.n150 OUT.t4 1191.28
R3994 OUT.n148 OUT.n147 1031.48
R3995 OUT.n149 OUT.n139 1031.48
R3996 OUT.n144 OUT.n143 963.661
R3997 OUT.n146 OUT.t3 948.736
R3998 OUT.n148 OUT.n140 877.239
R3999 OUT.t4 OUT.n149 877.239
R4000 OUT.n145 OUT.n141 854.746
R4001 OUT.n144 OUT.n142 841.893
R4002 OUT.n138 OUT.t1 222.722
R4003 OUT.n150 OUT.t5 207.718
R4004 OUT.n151 OUT.n68 185.824
R4005 OUT.n138 OUT.n137 163.862
R4006 OUT.n149 OUT.n148 154.24
R4007 OUT.n145 OUT.n144 137.116
R4008 OUT.n15 OUT.t2 64.755
R4009 OUT.n137 OUT.n102 49.503
R4010 OUT.n68 OUT.n33 49.503
R4011 OUT.n84 OUT.t0 42.441
R4012 OUT.n62 OUT.n61 32.833
R4013 OUT.n16 OUT.n15 30.553
R4014 OUT.n85 OUT.n84 29.289
R4015 OUT.n54 OUT.n53 26.863
R4016 OUT.n146 OUT.n145 24.1
R4017 OUT.n46 OUT.n45 20.893
R4018 OUT.n131 OUT.n130 20
R4019 OUT.n123 OUT.n122 16.363
R4020 OUT.n151 OUT.n150 15.198
R4021 OUT.n81 OUT.n80 15
R4022 OUT.n73 OUT.n72 15
R4023 OUT.n108 OUT.n107 15
R4024 OUT.n116 OUT.n115 15
R4025 OUT.n124 OUT.n123 15
R4026 OUT.n132 OUT.n131 15
R4027 OUT.n83 OUT.n82 15
R4028 OUT.n75 OUT.n74 15
R4029 OUT.n105 OUT.n104 15
R4030 OUT.n113 OUT.n112 15
R4031 OUT.n121 OUT.n120 15
R4032 OUT.n129 OUT.n128 15
R4033 OUT.n63 OUT.n62 15
R4034 OUT.n55 OUT.n54 15
R4035 OUT.n47 OUT.n46 15
R4036 OUT.n39 OUT.n38 15
R4037 OUT.n4 OUT.n3 15
R4038 OUT.n12 OUT.n11 15
R4039 OUT.n60 OUT.n59 15
R4040 OUT.n52 OUT.n51 15
R4041 OUT.n44 OUT.n43 15
R4042 OUT.n36 OUT.n35 15
R4043 OUT.n6 OUT.n5 15
R4044 OUT.n14 OUT.n13 15
R4045 OUT.n38 OUT.n37 14.924
R4046 OUT.n84 OUT.n83 14.586
R4047 OUT.n15 OUT.n14 14.123
R4048 OUT.n136 OUT.n135 13.634
R4049 OUT.n67 OUT.n66 13.544
R4050 OUT.n129 OUT.n127 12.917
R4051 OUT.n121 OUT.n119 12.917
R4052 OUT.n113 OUT.n111 12.917
R4053 OUT.n105 OUT.n103 12.917
R4054 OUT.n76 OUT.n75 12.917
R4055 OUT.n7 OUT.n6 12.917
R4056 OUT.n36 OUT.n34 12.917
R4057 OUT.n44 OUT.n42 12.917
R4058 OUT.n52 OUT.n50 12.917
R4059 OUT.n60 OUT.n58 12.917
R4060 OUT.n115 OUT.n114 12.727
R4061 OUT.n107 OUT.n106 9.09
R4062 OUT.n3 OUT.n2 8.954
R4063 OUT.n68 OUT.n67 8.805
R4064 OUT.n137 OUT.n136 8.695
R4065 OUT.n77 OUT.n76 5.741
R4066 OUT.n83 OUT.n81 5.741
R4067 OUT.n14 OUT.n12 5.741
R4068 OUT.n8 OUT.n7 5.741
R4069 OUT.n72 OUT.n71 5.454
R4070 OUT.n75 OUT.n73 5.023
R4071 OUT.n6 OUT.n4 5.023
R4072 OUT.n111 OUT.n110 4.305
R4073 OUT.n108 OUT.n105 4.305
R4074 OUT.n39 OUT.n36 4.305
R4075 OUT.n42 OUT.n41 4.305
R4076 OUT.n134 OUT.n133 3.947
R4077 OUT.n133 OUT.n132 3.947
R4078 OUT.n64 OUT.n63 3.947
R4079 OUT.n65 OUT.n64 3.947
R4080 OUT.n119 OUT.n118 3.588
R4081 OUT.n116 OUT.n113 3.588
R4082 OUT.n47 OUT.n44 3.588
R4083 OUT.n50 OUT.n49 3.588
R4084 OUT.n126 OUT.n125 3.229
R4085 OUT.n125 OUT.n124 3.229
R4086 OUT.n56 OUT.n55 3.229
R4087 OUT.n57 OUT.n56 3.229
R4088 OUT.n11 OUT.n10 2.984
R4089 OUT.n127 OUT.n126 2.87
R4090 OUT.n124 OUT.n121 2.87
R4091 OUT.n55 OUT.n52 2.87
R4092 OUT.n58 OUT.n57 2.87
R4093 OUT.n118 OUT.n117 2.511
R4094 OUT.n117 OUT.n116 2.511
R4095 OUT.n48 OUT.n47 2.511
R4096 OUT.n49 OUT.n48 2.511
R4097 OUT.n135 OUT.n134 2.152
R4098 OUT.n132 OUT.n129 2.152
R4099 OUT.n63 OUT.n60 2.152
R4100 OUT.n66 OUT.n65 2.152
R4101 OUT.n80 OUT.n79 1.818
R4102 OUT.n110 OUT.n109 1.794
R4103 OUT.n109 OUT.n108 1.794
R4104 OUT.n40 OUT.n39 1.794
R4105 OUT.n41 OUT.n40 1.794
R4106 OUT.n70 OUT.n69 1.076
R4107 OUT.n73 OUT.n70 1.076
R4108 OUT.n4 OUT.n1 1.076
R4109 OUT.n1 OUT.n0 1.076
R4110 OUT.n78 OUT.n77 0.358
R4111 OUT.n81 OUT.n78 0.358
R4112 OUT.n12 OUT.n9 0.358
R4113 OUT.n9 OUT.n8 0.358
R4114 OUT.n100 OUT.n99 0.144
R4115 OUT.n97 OUT.n96 0.144
R4116 OUT.n94 OUT.n93 0.144
R4117 OUT.n91 OUT.n90 0.144
R4118 OUT.n88 OUT.n87 0.144
R4119 OUT.n19 OUT.n18 0.144
R4120 OUT.n22 OUT.n21 0.144
R4121 OUT.n25 OUT.n24 0.144
R4122 OUT.n28 OUT.n27 0.144
R4123 OUT.n31 OUT.n30 0.144
R4124 OUT.n151 OUT.n138 0.129
R4125 OUT.n87 OUT.n86 0.043
R4126 OUT.n18 OUT.n17 0.043
R4127 OUT.n90 OUT.n89 0.038
R4128 OUT.n21 OUT.n20 0.038
R4129 OUT.n93 OUT.n92 0.032
R4130 OUT.n24 OUT.n23 0.032
R4131 OUT.n101 OUT.n100 0.029
R4132 OUT.n32 OUT.n31 0.029
R4133 OUT.n96 OUT.n95 0.027
R4134 OUT.n27 OUT.n26 0.027
R4135 OUT.n98 OUT.n97 0.024
R4136 OUT.n29 OUT.n28 0.024
R4137 OUT OUT.n151 0.022
R4138 OUT.n99 OUT.n98 0.021
R4139 OUT.n30 OUT.n29 0.021
R4140 OUT.n95 OUT.n94 0.019
R4141 OUT.n26 OUT.n25 0.019
R4142 OUT.n102 OUT.n101 0.016
R4143 OUT.n33 OUT.n32 0.016
R4144 OUT.n92 OUT.n91 0.013
R4145 OUT.n23 OUT.n22 0.013
R4146 OUT.n89 OUT.n88 0.008
R4147 OUT.n20 OUT.n19 0.008
R4148 OUT.n86 OUT.n85 0.002
R4149 OUT.n17 OUT.n16 0.002
R4150 a_1976_242.n96 a_1976_242.n95 1095.47
R4151 a_1976_242.n96 a_1976_242.n76 1093.38
R4152 a_1976_242.n97 a_1976_242.n57 1093.38
R4153 a_1976_242.n98 a_1976_242.n38 1093.36
R4154 a_1976_242.n19 a_1976_242.n18 1090.68
R4155 a_1976_242.n10 a_1976_242.n9 1025.05
R4156 a_1976_242.n2 a_1976_242.n1 1025.05
R4157 a_1976_242.n87 a_1976_242.n86 1025.05
R4158 a_1976_242.n79 a_1976_242.n78 1025.05
R4159 a_1976_242.n68 a_1976_242.n67 1025.05
R4160 a_1976_242.n59 a_1976_242.t5 1025.05
R4161 a_1976_242.n49 a_1976_242.t4 1025.05
R4162 a_1976_242.n41 a_1976_242.n40 1025.05
R4163 a_1976_242.n30 a_1976_242.t2 1025.05
R4164 a_1976_242.n22 a_1976_242.n21 1025.05
R4165 a_1976_242.n10 a_1976_242.n8 870.813
R4166 a_1976_242.n11 a_1976_242.n7 870.813
R4167 a_1976_242.n12 a_1976_242.n6 870.813
R4168 a_1976_242.n13 a_1976_242.t3 870.813
R4169 a_1976_242.n14 a_1976_242.n5 870.813
R4170 a_1976_242.n15 a_1976_242.n4 870.813
R4171 a_1976_242.n16 a_1976_242.n3 870.813
R4172 a_1976_242.n2 a_1976_242.n0 870.813
R4173 a_1976_242.n18 a_1976_242.n17 870.813
R4174 a_1976_242.n87 a_1976_242.t6 870.813
R4175 a_1976_242.n88 a_1976_242.n85 870.813
R4176 a_1976_242.n89 a_1976_242.n84 870.813
R4177 a_1976_242.n90 a_1976_242.n83 870.813
R4178 a_1976_242.n91 a_1976_242.n82 870.813
R4179 a_1976_242.n92 a_1976_242.n81 870.813
R4180 a_1976_242.n93 a_1976_242.n80 870.813
R4181 a_1976_242.n79 a_1976_242.n77 870.813
R4182 a_1976_242.n95 a_1976_242.n94 870.813
R4183 a_1976_242.n68 a_1976_242.n66 870.813
R4184 a_1976_242.n69 a_1976_242.n65 870.813
R4185 a_1976_242.n70 a_1976_242.n64 870.813
R4186 a_1976_242.n71 a_1976_242.n63 870.813
R4187 a_1976_242.n72 a_1976_242.n62 870.813
R4188 a_1976_242.n73 a_1976_242.n61 870.813
R4189 a_1976_242.n74 a_1976_242.n60 870.813
R4190 a_1976_242.n59 a_1976_242.n58 870.813
R4191 a_1976_242.n76 a_1976_242.n75 870.813
R4192 a_1976_242.n49 a_1976_242.n48 870.813
R4193 a_1976_242.n50 a_1976_242.n47 870.813
R4194 a_1976_242.n51 a_1976_242.n46 870.813
R4195 a_1976_242.n52 a_1976_242.n45 870.813
R4196 a_1976_242.n53 a_1976_242.n44 870.813
R4197 a_1976_242.n54 a_1976_242.n43 870.813
R4198 a_1976_242.n55 a_1976_242.n42 870.813
R4199 a_1976_242.n41 a_1976_242.n39 870.813
R4200 a_1976_242.n57 a_1976_242.n56 870.813
R4201 a_1976_242.n30 a_1976_242.n29 870.813
R4202 a_1976_242.n31 a_1976_242.n28 870.813
R4203 a_1976_242.n32 a_1976_242.n27 870.813
R4204 a_1976_242.n33 a_1976_242.n26 870.813
R4205 a_1976_242.n34 a_1976_242.n25 870.813
R4206 a_1976_242.n35 a_1976_242.n24 870.813
R4207 a_1976_242.n36 a_1976_242.n23 870.813
R4208 a_1976_242.n22 a_1976_242.n20 870.813
R4209 a_1976_242.n38 a_1976_242.n37 870.813
R4210 a_1976_242.t1 a_1976_242.n99 196.5
R4211 a_1976_242.n17 a_1976_242.n2 154.24
R4212 a_1976_242.n17 a_1976_242.n16 154.24
R4213 a_1976_242.n16 a_1976_242.n15 154.24
R4214 a_1976_242.n15 a_1976_242.n14 154.24
R4215 a_1976_242.n14 a_1976_242.n13 154.24
R4216 a_1976_242.n13 a_1976_242.n12 154.24
R4217 a_1976_242.n12 a_1976_242.n11 154.24
R4218 a_1976_242.n11 a_1976_242.n10 154.24
R4219 a_1976_242.n94 a_1976_242.n79 154.24
R4220 a_1976_242.n94 a_1976_242.n93 154.24
R4221 a_1976_242.n93 a_1976_242.n92 154.24
R4222 a_1976_242.n92 a_1976_242.n91 154.24
R4223 a_1976_242.n91 a_1976_242.n90 154.24
R4224 a_1976_242.n90 a_1976_242.n89 154.24
R4225 a_1976_242.n89 a_1976_242.n88 154.24
R4226 a_1976_242.n88 a_1976_242.n87 154.24
R4227 a_1976_242.n75 a_1976_242.n59 154.24
R4228 a_1976_242.n75 a_1976_242.n74 154.24
R4229 a_1976_242.n74 a_1976_242.n73 154.24
R4230 a_1976_242.n73 a_1976_242.n72 154.24
R4231 a_1976_242.n72 a_1976_242.n71 154.24
R4232 a_1976_242.n71 a_1976_242.n70 154.24
R4233 a_1976_242.n70 a_1976_242.n69 154.24
R4234 a_1976_242.n69 a_1976_242.n68 154.24
R4235 a_1976_242.n56 a_1976_242.n41 154.24
R4236 a_1976_242.n56 a_1976_242.n55 154.24
R4237 a_1976_242.n55 a_1976_242.n54 154.24
R4238 a_1976_242.n54 a_1976_242.n53 154.24
R4239 a_1976_242.n53 a_1976_242.n52 154.24
R4240 a_1976_242.n52 a_1976_242.n51 154.24
R4241 a_1976_242.n51 a_1976_242.n50 154.24
R4242 a_1976_242.n50 a_1976_242.n49 154.24
R4243 a_1976_242.n37 a_1976_242.n22 154.24
R4244 a_1976_242.n37 a_1976_242.n36 154.24
R4245 a_1976_242.n36 a_1976_242.n35 154.24
R4246 a_1976_242.n35 a_1976_242.n34 154.24
R4247 a_1976_242.n34 a_1976_242.n33 154.24
R4248 a_1976_242.n33 a_1976_242.n32 154.24
R4249 a_1976_242.n32 a_1976_242.n31 154.24
R4250 a_1976_242.n31 a_1976_242.n30 154.24
R4251 a_1976_242.n19 a_1976_242.t0 124.577
R4252 a_1976_242.n99 a_1976_242.n98 2.844
R4253 a_1976_242.n98 a_1976_242.n97 2.26
R4254 a_1976_242.n97 a_1976_242.n96 2.233
R4255 a_1976_242.n99 a_1976_242.n19 0.375
R4256 a_238_268.n174 a_238_268.n173 273.341
R4257 a_238_268.n184 a_238_268.n174 174.274
R4258 a_238_268.n174 a_238_268.n106 165.052
R4259 a_238_268.n106 a_238_268.n71 49.503
R4260 a_238_268.n173 a_238_268.n138 49.503
R4261 a_238_268.t2 a_238_268.n184 122.225
R4262 a_238_268.n55 a_238_268.t0 44.725
R4263 a_238_268.n122 a_238_268.t1 42.441
R4264 a_238_268.t2 a_238_268.n39 32.727
R4265 a_238_268.n56 a_238_268.n55 29.514
R4266 a_238_268.n123 a_238_268.n122 29.334
R4267 a_238_268.n39 a_238_268.n1 29.09
R4268 a_238_268.n100 a_238_268.n99 21.29
R4269 a_238_268.n167 a_238_268.n166 20
R4270 a_238_268.n178 a_238_268.n177 20
R4271 a_238_268.n92 a_238_268.n91 17.419
R4272 a_238_268.n159 a_238_268.n158 16.363
R4273 a_238_268.n6 a_238_268.n5 16.363
R4274 a_238_268.n101 a_238_268.n100 15
R4275 a_238_268.n93 a_238_268.n92 15
R4276 a_238_268.n85 a_238_268.n84 15
R4277 a_238_268.n77 a_238_268.n76 15
R4278 a_238_268.n44 a_238_268.n43 15
R4279 a_238_268.n52 a_238_268.n51 15
R4280 a_238_268.n98 a_238_268.n97 15
R4281 a_238_268.n90 a_238_268.n89 15
R4282 a_238_268.n82 a_238_268.n81 15
R4283 a_238_268.n74 a_238_268.n73 15
R4284 a_238_268.n46 a_238_268.n45 15
R4285 a_238_268.n54 a_238_268.n53 15
R4286 a_238_268.n119 a_238_268.n118 15
R4287 a_238_268.n111 a_238_268.n110 15
R4288 a_238_268.n144 a_238_268.n143 15
R4289 a_238_268.n152 a_238_268.n151 15
R4290 a_238_268.n160 a_238_268.n159 15
R4291 a_238_268.n168 a_238_268.n167 15
R4292 a_238_268.n121 a_238_268.n120 15
R4293 a_238_268.n113 a_238_268.n112 15
R4294 a_238_268.n141 a_238_268.n140 15
R4295 a_238_268.n149 a_238_268.n148 15
R4296 a_238_268.n157 a_238_268.n156 15
R4297 a_238_268.n165 a_238_268.n164 15
R4298 a_238_268.n31 a_238_268.n30 15
R4299 a_238_268.n23 a_238_268.n22 15
R4300 a_238_268.n15 a_238_268.n14 15
R4301 a_238_268.n7 a_238_268.n6 15
R4302 a_238_268.n179 a_238_268.n178 15
R4303 a_238_268.n39 a_238_268.n38 15
R4304 a_238_268.n33 a_238_268.n32 15
R4305 a_238_268.n25 a_238_268.n24 15
R4306 a_238_268.n17 a_238_268.n16 15
R4307 a_238_268.n9 a_238_268.n8 15
R4308 a_238_268.n176 a_238_268.n175 15
R4309 a_238_268.n122 a_238_268.n121 14.586
R4310 a_238_268.n55 a_238_268.n54 14.523
R4311 a_238_268.n172 a_238_268.n171 13.634
R4312 a_238_268.n183 a_238_268.n182 13.634
R4313 a_238_268.n105 a_238_268.n104 13.624
R4314 a_238_268.n84 a_238_268.n83 13.548
R4315 a_238_268.n47 a_238_268.n46 12.917
R4316 a_238_268.n74 a_238_268.n72 12.917
R4317 a_238_268.n82 a_238_268.n80 12.917
R4318 a_238_268.n90 a_238_268.n88 12.917
R4319 a_238_268.n98 a_238_268.n96 12.917
R4320 a_238_268.n165 a_238_268.n163 12.917
R4321 a_238_268.n157 a_238_268.n155 12.917
R4322 a_238_268.n149 a_238_268.n147 12.917
R4323 a_238_268.n141 a_238_268.n139 12.917
R4324 a_238_268.n114 a_238_268.n113 12.917
R4325 a_238_268.n10 a_238_268.n9 12.917
R4326 a_238_268.n18 a_238_268.n17 12.917
R4327 a_238_268.n26 a_238_268.n25 12.917
R4328 a_238_268.n34 a_238_268.n33 12.917
R4329 a_238_268.n151 a_238_268.n150 12.727
R4330 a_238_268.n14 a_238_268.n13 12.727
R4331 a_238_268.n76 a_238_268.n75 9.677
R4332 a_238_268.n143 a_238_268.n142 9.09
R4333 a_238_268.n22 a_238_268.n21 9.09
R4334 a_238_268.n106 a_238_268.n105 8.708
R4335 a_238_268.n173 a_238_268.n172 8.695
R4336 a_238_268.n184 a_238_268.n183 8.695
R4337 a_238_268.n43 a_238_268.n42 5.806
R4338 a_238_268.n54 a_238_268.n52 5.741
R4339 a_238_268.n48 a_238_268.n47 5.741
R4340 a_238_268.n115 a_238_268.n114 5.741
R4341 a_238_268.n121 a_238_268.n119 5.741
R4342 a_238_268.n35 a_238_268.n34 5.741
R4343 a_238_268.n38 a_238_268.n37 5.741
R4344 a_238_268.n110 a_238_268.n109 5.454
R4345 a_238_268.n30 a_238_268.n29 5.454
R4346 a_238_268.n46 a_238_268.n44 5.023
R4347 a_238_268.n113 a_238_268.n111 5.023
R4348 a_238_268.n27 a_238_268.n26 5.023
R4349 a_238_268.n33 a_238_268.n31 5.023
R4350 a_238_268.n77 a_238_268.n74 4.305
R4351 a_238_268.n80 a_238_268.n79 4.305
R4352 a_238_268.n147 a_238_268.n146 4.305
R4353 a_238_268.n144 a_238_268.n141 4.305
R4354 a_238_268.n19 a_238_268.n18 4.305
R4355 a_238_268.n25 a_238_268.n23 4.305
R4356 a_238_268.n102 a_238_268.n101 3.947
R4357 a_238_268.n103 a_238_268.n102 3.947
R4358 a_238_268.n170 a_238_268.n169 3.947
R4359 a_238_268.n169 a_238_268.n168 3.947
R4360 a_238_268.n181 a_238_268.n180 3.947
R4361 a_238_268.n180 a_238_268.n179 3.947
R4362 a_238_268.n85 a_238_268.n82 3.588
R4363 a_238_268.n88 a_238_268.n87 3.588
R4364 a_238_268.n155 a_238_268.n154 3.588
R4365 a_238_268.n152 a_238_268.n149 3.588
R4366 a_238_268.n11 a_238_268.n10 3.588
R4367 a_238_268.n17 a_238_268.n15 3.588
R4368 a_238_268.n94 a_238_268.n93 3.229
R4369 a_238_268.n95 a_238_268.n94 3.229
R4370 a_238_268.n162 a_238_268.n161 3.229
R4371 a_238_268.n161 a_238_268.n160 3.229
R4372 a_238_268.n4 a_238_268.n3 3.229
R4373 a_238_268.n7 a_238_268.n4 3.229
R4374 a_238_268.n93 a_238_268.n90 2.87
R4375 a_238_268.n96 a_238_268.n95 2.87
R4376 a_238_268.n163 a_238_268.n162 2.87
R4377 a_238_268.n160 a_238_268.n157 2.87
R4378 a_238_268.n3 a_238_268.n2 2.87
R4379 a_238_268.n9 a_238_268.n7 2.87
R4380 a_238_268.n86 a_238_268.n85 2.511
R4381 a_238_268.n87 a_238_268.n86 2.511
R4382 a_238_268.n154 a_238_268.n153 2.511
R4383 a_238_268.n153 a_238_268.n152 2.511
R4384 a_238_268.n12 a_238_268.n11 2.511
R4385 a_238_268.n15 a_238_268.n12 2.511
R4386 a_238_268.n101 a_238_268.n98 2.152
R4387 a_238_268.n104 a_238_268.n103 2.152
R4388 a_238_268.n171 a_238_268.n170 2.152
R4389 a_238_268.n168 a_238_268.n165 2.152
R4390 a_238_268.n182 a_238_268.n181 2.152
R4391 a_238_268.n179 a_238_268.n176 2.152
R4392 a_238_268.n51 a_238_268.n50 1.935
R4393 a_238_268.n118 a_238_268.n117 1.818
R4394 a_238_268.n1 a_238_268.n0 1.818
R4395 a_238_268.n78 a_238_268.n77 1.794
R4396 a_238_268.n79 a_238_268.n78 1.794
R4397 a_238_268.n146 a_238_268.n145 1.794
R4398 a_238_268.n145 a_238_268.n144 1.794
R4399 a_238_268.n20 a_238_268.n19 1.794
R4400 a_238_268.n23 a_238_268.n20 1.794
R4401 a_238_268.n44 a_238_268.n41 1.076
R4402 a_238_268.n41 a_238_268.n40 1.076
R4403 a_238_268.n108 a_238_268.n107 1.076
R4404 a_238_268.n111 a_238_268.n108 1.076
R4405 a_238_268.n28 a_238_268.n27 1.076
R4406 a_238_268.n31 a_238_268.n28 1.076
R4407 a_238_268.n52 a_238_268.n49 0.358
R4408 a_238_268.n49 a_238_268.n48 0.358
R4409 a_238_268.n116 a_238_268.n115 0.358
R4410 a_238_268.n119 a_238_268.n116 0.358
R4411 a_238_268.n36 a_238_268.n35 0.358
R4412 a_238_268.n37 a_238_268.n36 0.358
R4413 a_238_268.n57 a_238_268.n56 0.144
R4414 a_238_268.n60 a_238_268.n59 0.144
R4415 a_238_268.n63 a_238_268.n62 0.144
R4416 a_238_268.n66 a_238_268.n65 0.144
R4417 a_238_268.n69 a_238_268.n68 0.144
R4418 a_238_268.n136 a_238_268.n135 0.144
R4419 a_238_268.n133 a_238_268.n132 0.144
R4420 a_238_268.n130 a_238_268.n129 0.144
R4421 a_238_268.n127 a_238_268.n126 0.144
R4422 a_238_268.n124 a_238_268.n123 0.144
R4423 a_238_268.n59 a_238_268.n58 0.038
R4424 a_238_268.n126 a_238_268.n125 0.038
R4425 a_238_268.n62 a_238_268.n61 0.032
R4426 a_238_268.n129 a_238_268.n128 0.032
R4427 a_238_268.n70 a_238_268.n69 0.029
R4428 a_238_268.n137 a_238_268.n136 0.029
R4429 a_238_268.n65 a_238_268.n64 0.027
R4430 a_238_268.n132 a_238_268.n131 0.027
R4431 a_238_268.n67 a_238_268.n66 0.024
R4432 a_238_268.n134 a_238_268.n133 0.024
R4433 a_238_268.n68 a_238_268.n67 0.021
R4434 a_238_268.n135 a_238_268.n134 0.021
R4435 a_238_268.n64 a_238_268.n63 0.019
R4436 a_238_268.n131 a_238_268.n130 0.019
R4437 a_238_268.n71 a_238_268.n70 0.016
R4438 a_238_268.n138 a_238_268.n137 0.016
R4439 a_238_268.n61 a_238_268.n60 0.013
R4440 a_238_268.n128 a_238_268.n127 0.013
R4441 a_238_268.n58 a_238_268.n57 0.008
R4442 a_238_268.n125 a_238_268.n124 0.008
R4443 a_12468_224.n184 a_12468_224.n174 312.09
R4444 a_12468_224.n174 a_12468_224.n106 165.03
R4445 a_12468_224.n174 a_12468_224.n173 139.83
R4446 a_12468_224.n106 a_12468_224.n71 49.503
R4447 a_12468_224.n173 a_12468_224.n138 49.503
R4448 a_12468_224.t2 a_12468_224.n184 122.225
R4449 a_12468_224.n55 a_12468_224.t0 44.725
R4450 a_12468_224.n122 a_12468_224.t1 42.441
R4451 a_12468_224.t2 a_12468_224.n39 32.727
R4452 a_12468_224.n56 a_12468_224.n55 29.514
R4453 a_12468_224.n123 a_12468_224.n122 29.334
R4454 a_12468_224.n39 a_12468_224.n1 29.09
R4455 a_12468_224.n100 a_12468_224.n99 21.29
R4456 a_12468_224.n167 a_12468_224.n166 20
R4457 a_12468_224.n178 a_12468_224.n177 20
R4458 a_12468_224.n92 a_12468_224.n91 17.419
R4459 a_12468_224.n159 a_12468_224.n158 16.363
R4460 a_12468_224.n6 a_12468_224.n5 16.363
R4461 a_12468_224.n101 a_12468_224.n100 15
R4462 a_12468_224.n93 a_12468_224.n92 15
R4463 a_12468_224.n85 a_12468_224.n84 15
R4464 a_12468_224.n77 a_12468_224.n76 15
R4465 a_12468_224.n44 a_12468_224.n43 15
R4466 a_12468_224.n52 a_12468_224.n51 15
R4467 a_12468_224.n98 a_12468_224.n97 15
R4468 a_12468_224.n90 a_12468_224.n89 15
R4469 a_12468_224.n82 a_12468_224.n81 15
R4470 a_12468_224.n74 a_12468_224.n73 15
R4471 a_12468_224.n46 a_12468_224.n45 15
R4472 a_12468_224.n54 a_12468_224.n53 15
R4473 a_12468_224.n119 a_12468_224.n118 15
R4474 a_12468_224.n111 a_12468_224.n110 15
R4475 a_12468_224.n144 a_12468_224.n143 15
R4476 a_12468_224.n152 a_12468_224.n151 15
R4477 a_12468_224.n160 a_12468_224.n159 15
R4478 a_12468_224.n168 a_12468_224.n167 15
R4479 a_12468_224.n121 a_12468_224.n120 15
R4480 a_12468_224.n113 a_12468_224.n112 15
R4481 a_12468_224.n141 a_12468_224.n140 15
R4482 a_12468_224.n149 a_12468_224.n148 15
R4483 a_12468_224.n157 a_12468_224.n156 15
R4484 a_12468_224.n165 a_12468_224.n164 15
R4485 a_12468_224.n31 a_12468_224.n30 15
R4486 a_12468_224.n23 a_12468_224.n22 15
R4487 a_12468_224.n15 a_12468_224.n14 15
R4488 a_12468_224.n7 a_12468_224.n6 15
R4489 a_12468_224.n179 a_12468_224.n178 15
R4490 a_12468_224.n39 a_12468_224.n38 15
R4491 a_12468_224.n33 a_12468_224.n32 15
R4492 a_12468_224.n25 a_12468_224.n24 15
R4493 a_12468_224.n17 a_12468_224.n16 15
R4494 a_12468_224.n9 a_12468_224.n8 15
R4495 a_12468_224.n176 a_12468_224.n175 15
R4496 a_12468_224.n122 a_12468_224.n121 14.586
R4497 a_12468_224.n55 a_12468_224.n54 14.523
R4498 a_12468_224.n172 a_12468_224.n171 13.634
R4499 a_12468_224.n183 a_12468_224.n182 13.634
R4500 a_12468_224.n105 a_12468_224.n104 13.624
R4501 a_12468_224.n84 a_12468_224.n83 13.548
R4502 a_12468_224.n47 a_12468_224.n46 12.917
R4503 a_12468_224.n74 a_12468_224.n72 12.917
R4504 a_12468_224.n82 a_12468_224.n80 12.917
R4505 a_12468_224.n90 a_12468_224.n88 12.917
R4506 a_12468_224.n98 a_12468_224.n96 12.917
R4507 a_12468_224.n165 a_12468_224.n163 12.917
R4508 a_12468_224.n157 a_12468_224.n155 12.917
R4509 a_12468_224.n149 a_12468_224.n147 12.917
R4510 a_12468_224.n141 a_12468_224.n139 12.917
R4511 a_12468_224.n114 a_12468_224.n113 12.917
R4512 a_12468_224.n10 a_12468_224.n9 12.917
R4513 a_12468_224.n18 a_12468_224.n17 12.917
R4514 a_12468_224.n26 a_12468_224.n25 12.917
R4515 a_12468_224.n34 a_12468_224.n33 12.917
R4516 a_12468_224.n151 a_12468_224.n150 12.727
R4517 a_12468_224.n14 a_12468_224.n13 12.727
R4518 a_12468_224.n76 a_12468_224.n75 9.677
R4519 a_12468_224.n143 a_12468_224.n142 9.09
R4520 a_12468_224.n22 a_12468_224.n21 9.09
R4521 a_12468_224.n106 a_12468_224.n105 8.708
R4522 a_12468_224.n173 a_12468_224.n172 8.695
R4523 a_12468_224.n184 a_12468_224.n183 8.695
R4524 a_12468_224.n43 a_12468_224.n42 5.806
R4525 a_12468_224.n54 a_12468_224.n52 5.741
R4526 a_12468_224.n48 a_12468_224.n47 5.741
R4527 a_12468_224.n115 a_12468_224.n114 5.741
R4528 a_12468_224.n121 a_12468_224.n119 5.741
R4529 a_12468_224.n35 a_12468_224.n34 5.741
R4530 a_12468_224.n38 a_12468_224.n37 5.741
R4531 a_12468_224.n110 a_12468_224.n109 5.454
R4532 a_12468_224.n30 a_12468_224.n29 5.454
R4533 a_12468_224.n46 a_12468_224.n44 5.023
R4534 a_12468_224.n113 a_12468_224.n111 5.023
R4535 a_12468_224.n27 a_12468_224.n26 5.023
R4536 a_12468_224.n33 a_12468_224.n31 5.023
R4537 a_12468_224.n77 a_12468_224.n74 4.305
R4538 a_12468_224.n80 a_12468_224.n79 4.305
R4539 a_12468_224.n147 a_12468_224.n146 4.305
R4540 a_12468_224.n144 a_12468_224.n141 4.305
R4541 a_12468_224.n19 a_12468_224.n18 4.305
R4542 a_12468_224.n25 a_12468_224.n23 4.305
R4543 a_12468_224.n102 a_12468_224.n101 3.947
R4544 a_12468_224.n103 a_12468_224.n102 3.947
R4545 a_12468_224.n170 a_12468_224.n169 3.947
R4546 a_12468_224.n169 a_12468_224.n168 3.947
R4547 a_12468_224.n181 a_12468_224.n180 3.947
R4548 a_12468_224.n180 a_12468_224.n179 3.947
R4549 a_12468_224.n85 a_12468_224.n82 3.588
R4550 a_12468_224.n88 a_12468_224.n87 3.588
R4551 a_12468_224.n155 a_12468_224.n154 3.588
R4552 a_12468_224.n152 a_12468_224.n149 3.588
R4553 a_12468_224.n11 a_12468_224.n10 3.588
R4554 a_12468_224.n17 a_12468_224.n15 3.588
R4555 a_12468_224.n94 a_12468_224.n93 3.229
R4556 a_12468_224.n95 a_12468_224.n94 3.229
R4557 a_12468_224.n162 a_12468_224.n161 3.229
R4558 a_12468_224.n161 a_12468_224.n160 3.229
R4559 a_12468_224.n4 a_12468_224.n3 3.229
R4560 a_12468_224.n7 a_12468_224.n4 3.229
R4561 a_12468_224.n93 a_12468_224.n90 2.87
R4562 a_12468_224.n96 a_12468_224.n95 2.87
R4563 a_12468_224.n163 a_12468_224.n162 2.87
R4564 a_12468_224.n160 a_12468_224.n157 2.87
R4565 a_12468_224.n3 a_12468_224.n2 2.87
R4566 a_12468_224.n9 a_12468_224.n7 2.87
R4567 a_12468_224.n86 a_12468_224.n85 2.511
R4568 a_12468_224.n87 a_12468_224.n86 2.511
R4569 a_12468_224.n154 a_12468_224.n153 2.511
R4570 a_12468_224.n153 a_12468_224.n152 2.511
R4571 a_12468_224.n12 a_12468_224.n11 2.511
R4572 a_12468_224.n15 a_12468_224.n12 2.511
R4573 a_12468_224.n101 a_12468_224.n98 2.152
R4574 a_12468_224.n104 a_12468_224.n103 2.152
R4575 a_12468_224.n171 a_12468_224.n170 2.152
R4576 a_12468_224.n168 a_12468_224.n165 2.152
R4577 a_12468_224.n182 a_12468_224.n181 2.152
R4578 a_12468_224.n179 a_12468_224.n176 2.152
R4579 a_12468_224.n51 a_12468_224.n50 1.935
R4580 a_12468_224.n118 a_12468_224.n117 1.818
R4581 a_12468_224.n1 a_12468_224.n0 1.818
R4582 a_12468_224.n78 a_12468_224.n77 1.794
R4583 a_12468_224.n79 a_12468_224.n78 1.794
R4584 a_12468_224.n146 a_12468_224.n145 1.794
R4585 a_12468_224.n145 a_12468_224.n144 1.794
R4586 a_12468_224.n20 a_12468_224.n19 1.794
R4587 a_12468_224.n23 a_12468_224.n20 1.794
R4588 a_12468_224.n44 a_12468_224.n41 1.076
R4589 a_12468_224.n41 a_12468_224.n40 1.076
R4590 a_12468_224.n108 a_12468_224.n107 1.076
R4591 a_12468_224.n111 a_12468_224.n108 1.076
R4592 a_12468_224.n28 a_12468_224.n27 1.076
R4593 a_12468_224.n31 a_12468_224.n28 1.076
R4594 a_12468_224.n52 a_12468_224.n49 0.358
R4595 a_12468_224.n49 a_12468_224.n48 0.358
R4596 a_12468_224.n116 a_12468_224.n115 0.358
R4597 a_12468_224.n119 a_12468_224.n116 0.358
R4598 a_12468_224.n36 a_12468_224.n35 0.358
R4599 a_12468_224.n37 a_12468_224.n36 0.358
R4600 a_12468_224.n57 a_12468_224.n56 0.144
R4601 a_12468_224.n60 a_12468_224.n59 0.144
R4602 a_12468_224.n63 a_12468_224.n62 0.144
R4603 a_12468_224.n66 a_12468_224.n65 0.144
R4604 a_12468_224.n69 a_12468_224.n68 0.144
R4605 a_12468_224.n136 a_12468_224.n135 0.144
R4606 a_12468_224.n133 a_12468_224.n132 0.144
R4607 a_12468_224.n130 a_12468_224.n129 0.144
R4608 a_12468_224.n127 a_12468_224.n126 0.144
R4609 a_12468_224.n124 a_12468_224.n123 0.144
R4610 a_12468_224.n59 a_12468_224.n58 0.038
R4611 a_12468_224.n126 a_12468_224.n125 0.038
R4612 a_12468_224.n62 a_12468_224.n61 0.032
R4613 a_12468_224.n129 a_12468_224.n128 0.032
R4614 a_12468_224.n70 a_12468_224.n69 0.029
R4615 a_12468_224.n137 a_12468_224.n136 0.029
R4616 a_12468_224.n65 a_12468_224.n64 0.027
R4617 a_12468_224.n132 a_12468_224.n131 0.027
R4618 a_12468_224.n67 a_12468_224.n66 0.024
R4619 a_12468_224.n134 a_12468_224.n133 0.024
R4620 a_12468_224.n68 a_12468_224.n67 0.021
R4621 a_12468_224.n135 a_12468_224.n134 0.021
R4622 a_12468_224.n64 a_12468_224.n63 0.019
R4623 a_12468_224.n131 a_12468_224.n130 0.019
R4624 a_12468_224.n71 a_12468_224.n70 0.016
R4625 a_12468_224.n138 a_12468_224.n137 0.016
R4626 a_12468_224.n61 a_12468_224.n60 0.013
R4627 a_12468_224.n128 a_12468_224.n127 0.013
R4628 a_12468_224.n58 a_12468_224.n57 0.008
R4629 a_12468_224.n125 a_12468_224.n124 0.008
R4630 a_6224_252.n184 a_6224_252.n174 312.007
R4631 a_6224_252.n174 a_6224_252.n173 273.226
R4632 a_6224_252.n174 a_6224_252.n106 165.052
R4633 a_6224_252.n106 a_6224_252.n71 49.503
R4634 a_6224_252.n173 a_6224_252.n138 49.503
R4635 a_6224_252.t1 a_6224_252.n184 122.225
R4636 a_6224_252.n55 a_6224_252.t2 42.441
R4637 a_6224_252.n122 a_6224_252.t0 42.441
R4638 a_6224_252.t1 a_6224_252.n39 32.727
R4639 a_6224_252.n56 a_6224_252.n55 29.334
R4640 a_6224_252.n123 a_6224_252.n122 29.334
R4641 a_6224_252.n39 a_6224_252.n1 29.09
R4642 a_6224_252.n100 a_6224_252.n99 20
R4643 a_6224_252.n167 a_6224_252.n166 20
R4644 a_6224_252.n178 a_6224_252.n177 20
R4645 a_6224_252.n92 a_6224_252.n91 16.363
R4646 a_6224_252.n159 a_6224_252.n158 16.363
R4647 a_6224_252.n6 a_6224_252.n5 16.363
R4648 a_6224_252.n52 a_6224_252.n51 15
R4649 a_6224_252.n44 a_6224_252.n43 15
R4650 a_6224_252.n77 a_6224_252.n76 15
R4651 a_6224_252.n85 a_6224_252.n84 15
R4652 a_6224_252.n93 a_6224_252.n92 15
R4653 a_6224_252.n54 a_6224_252.n53 15
R4654 a_6224_252.n46 a_6224_252.n45 15
R4655 a_6224_252.n74 a_6224_252.n73 15
R4656 a_6224_252.n82 a_6224_252.n81 15
R4657 a_6224_252.n90 a_6224_252.n89 15
R4658 a_6224_252.n98 a_6224_252.n97 15
R4659 a_6224_252.n101 a_6224_252.n100 15
R4660 a_6224_252.n119 a_6224_252.n118 15
R4661 a_6224_252.n111 a_6224_252.n110 15
R4662 a_6224_252.n144 a_6224_252.n143 15
R4663 a_6224_252.n152 a_6224_252.n151 15
R4664 a_6224_252.n160 a_6224_252.n159 15
R4665 a_6224_252.n168 a_6224_252.n167 15
R4666 a_6224_252.n121 a_6224_252.n120 15
R4667 a_6224_252.n113 a_6224_252.n112 15
R4668 a_6224_252.n141 a_6224_252.n140 15
R4669 a_6224_252.n149 a_6224_252.n148 15
R4670 a_6224_252.n157 a_6224_252.n156 15
R4671 a_6224_252.n165 a_6224_252.n164 15
R4672 a_6224_252.n31 a_6224_252.n30 15
R4673 a_6224_252.n23 a_6224_252.n22 15
R4674 a_6224_252.n15 a_6224_252.n14 15
R4675 a_6224_252.n7 a_6224_252.n6 15
R4676 a_6224_252.n179 a_6224_252.n178 15
R4677 a_6224_252.n39 a_6224_252.n38 15
R4678 a_6224_252.n33 a_6224_252.n32 15
R4679 a_6224_252.n25 a_6224_252.n24 15
R4680 a_6224_252.n17 a_6224_252.n16 15
R4681 a_6224_252.n9 a_6224_252.n8 15
R4682 a_6224_252.n176 a_6224_252.n175 15
R4683 a_6224_252.n55 a_6224_252.n54 14.586
R4684 a_6224_252.n122 a_6224_252.n121 14.586
R4685 a_6224_252.n105 a_6224_252.n104 13.634
R4686 a_6224_252.n172 a_6224_252.n171 13.634
R4687 a_6224_252.n183 a_6224_252.n182 13.634
R4688 a_6224_252.n47 a_6224_252.n46 12.917
R4689 a_6224_252.n74 a_6224_252.n72 12.917
R4690 a_6224_252.n82 a_6224_252.n80 12.917
R4691 a_6224_252.n90 a_6224_252.n88 12.917
R4692 a_6224_252.n98 a_6224_252.n96 12.917
R4693 a_6224_252.n165 a_6224_252.n163 12.917
R4694 a_6224_252.n157 a_6224_252.n155 12.917
R4695 a_6224_252.n149 a_6224_252.n147 12.917
R4696 a_6224_252.n141 a_6224_252.n139 12.917
R4697 a_6224_252.n114 a_6224_252.n113 12.917
R4698 a_6224_252.n10 a_6224_252.n9 12.917
R4699 a_6224_252.n18 a_6224_252.n17 12.917
R4700 a_6224_252.n26 a_6224_252.n25 12.917
R4701 a_6224_252.n34 a_6224_252.n33 12.917
R4702 a_6224_252.n84 a_6224_252.n83 12.727
R4703 a_6224_252.n151 a_6224_252.n150 12.727
R4704 a_6224_252.n14 a_6224_252.n13 12.727
R4705 a_6224_252.n76 a_6224_252.n75 9.09
R4706 a_6224_252.n143 a_6224_252.n142 9.09
R4707 a_6224_252.n22 a_6224_252.n21 9.09
R4708 a_6224_252.n106 a_6224_252.n105 8.695
R4709 a_6224_252.n173 a_6224_252.n172 8.695
R4710 a_6224_252.n184 a_6224_252.n183 8.695
R4711 a_6224_252.n54 a_6224_252.n52 5.741
R4712 a_6224_252.n48 a_6224_252.n47 5.741
R4713 a_6224_252.n115 a_6224_252.n114 5.741
R4714 a_6224_252.n121 a_6224_252.n119 5.741
R4715 a_6224_252.n35 a_6224_252.n34 5.741
R4716 a_6224_252.n38 a_6224_252.n37 5.741
R4717 a_6224_252.n43 a_6224_252.n42 5.454
R4718 a_6224_252.n110 a_6224_252.n109 5.454
R4719 a_6224_252.n30 a_6224_252.n29 5.454
R4720 a_6224_252.n46 a_6224_252.n44 5.023
R4721 a_6224_252.n113 a_6224_252.n111 5.023
R4722 a_6224_252.n27 a_6224_252.n26 5.023
R4723 a_6224_252.n33 a_6224_252.n31 5.023
R4724 a_6224_252.n77 a_6224_252.n74 4.305
R4725 a_6224_252.n80 a_6224_252.n79 4.305
R4726 a_6224_252.n147 a_6224_252.n146 4.305
R4727 a_6224_252.n144 a_6224_252.n141 4.305
R4728 a_6224_252.n19 a_6224_252.n18 4.305
R4729 a_6224_252.n25 a_6224_252.n23 4.305
R4730 a_6224_252.n102 a_6224_252.n101 3.947
R4731 a_6224_252.n103 a_6224_252.n102 3.947
R4732 a_6224_252.n170 a_6224_252.n169 3.947
R4733 a_6224_252.n169 a_6224_252.n168 3.947
R4734 a_6224_252.n181 a_6224_252.n180 3.947
R4735 a_6224_252.n180 a_6224_252.n179 3.947
R4736 a_6224_252.n85 a_6224_252.n82 3.588
R4737 a_6224_252.n88 a_6224_252.n87 3.588
R4738 a_6224_252.n155 a_6224_252.n154 3.588
R4739 a_6224_252.n152 a_6224_252.n149 3.588
R4740 a_6224_252.n11 a_6224_252.n10 3.588
R4741 a_6224_252.n17 a_6224_252.n15 3.588
R4742 a_6224_252.n94 a_6224_252.n93 3.229
R4743 a_6224_252.n95 a_6224_252.n94 3.229
R4744 a_6224_252.n162 a_6224_252.n161 3.229
R4745 a_6224_252.n161 a_6224_252.n160 3.229
R4746 a_6224_252.n4 a_6224_252.n3 3.229
R4747 a_6224_252.n7 a_6224_252.n4 3.229
R4748 a_6224_252.n93 a_6224_252.n90 2.87
R4749 a_6224_252.n96 a_6224_252.n95 2.87
R4750 a_6224_252.n163 a_6224_252.n162 2.87
R4751 a_6224_252.n160 a_6224_252.n157 2.87
R4752 a_6224_252.n3 a_6224_252.n2 2.87
R4753 a_6224_252.n9 a_6224_252.n7 2.87
R4754 a_6224_252.n86 a_6224_252.n85 2.511
R4755 a_6224_252.n87 a_6224_252.n86 2.511
R4756 a_6224_252.n154 a_6224_252.n153 2.511
R4757 a_6224_252.n153 a_6224_252.n152 2.511
R4758 a_6224_252.n12 a_6224_252.n11 2.511
R4759 a_6224_252.n15 a_6224_252.n12 2.511
R4760 a_6224_252.n101 a_6224_252.n98 2.152
R4761 a_6224_252.n104 a_6224_252.n103 2.152
R4762 a_6224_252.n171 a_6224_252.n170 2.152
R4763 a_6224_252.n168 a_6224_252.n165 2.152
R4764 a_6224_252.n182 a_6224_252.n181 2.152
R4765 a_6224_252.n179 a_6224_252.n176 2.152
R4766 a_6224_252.n51 a_6224_252.n50 1.818
R4767 a_6224_252.n118 a_6224_252.n117 1.818
R4768 a_6224_252.n1 a_6224_252.n0 1.818
R4769 a_6224_252.n78 a_6224_252.n77 1.794
R4770 a_6224_252.n79 a_6224_252.n78 1.794
R4771 a_6224_252.n146 a_6224_252.n145 1.794
R4772 a_6224_252.n145 a_6224_252.n144 1.794
R4773 a_6224_252.n20 a_6224_252.n19 1.794
R4774 a_6224_252.n23 a_6224_252.n20 1.794
R4775 a_6224_252.n44 a_6224_252.n41 1.076
R4776 a_6224_252.n41 a_6224_252.n40 1.076
R4777 a_6224_252.n108 a_6224_252.n107 1.076
R4778 a_6224_252.n111 a_6224_252.n108 1.076
R4779 a_6224_252.n28 a_6224_252.n27 1.076
R4780 a_6224_252.n31 a_6224_252.n28 1.076
R4781 a_6224_252.n52 a_6224_252.n49 0.358
R4782 a_6224_252.n49 a_6224_252.n48 0.358
R4783 a_6224_252.n116 a_6224_252.n115 0.358
R4784 a_6224_252.n119 a_6224_252.n116 0.358
R4785 a_6224_252.n36 a_6224_252.n35 0.358
R4786 a_6224_252.n37 a_6224_252.n36 0.358
R4787 a_6224_252.n57 a_6224_252.n56 0.144
R4788 a_6224_252.n60 a_6224_252.n59 0.144
R4789 a_6224_252.n63 a_6224_252.n62 0.144
R4790 a_6224_252.n66 a_6224_252.n65 0.144
R4791 a_6224_252.n69 a_6224_252.n68 0.144
R4792 a_6224_252.n136 a_6224_252.n135 0.144
R4793 a_6224_252.n133 a_6224_252.n132 0.144
R4794 a_6224_252.n130 a_6224_252.n129 0.144
R4795 a_6224_252.n127 a_6224_252.n126 0.144
R4796 a_6224_252.n124 a_6224_252.n123 0.144
R4797 a_6224_252.n59 a_6224_252.n58 0.038
R4798 a_6224_252.n126 a_6224_252.n125 0.038
R4799 a_6224_252.n62 a_6224_252.n61 0.032
R4800 a_6224_252.n129 a_6224_252.n128 0.032
R4801 a_6224_252.n70 a_6224_252.n69 0.029
R4802 a_6224_252.n137 a_6224_252.n136 0.029
R4803 a_6224_252.n65 a_6224_252.n64 0.027
R4804 a_6224_252.n132 a_6224_252.n131 0.027
R4805 a_6224_252.n67 a_6224_252.n66 0.024
R4806 a_6224_252.n134 a_6224_252.n133 0.024
R4807 a_6224_252.n68 a_6224_252.n67 0.021
R4808 a_6224_252.n135 a_6224_252.n134 0.021
R4809 a_6224_252.n64 a_6224_252.n63 0.019
R4810 a_6224_252.n131 a_6224_252.n130 0.019
R4811 a_6224_252.n71 a_6224_252.n70 0.016
R4812 a_6224_252.n138 a_6224_252.n137 0.016
R4813 a_6224_252.n61 a_6224_252.n60 0.013
R4814 a_6224_252.n128 a_6224_252.n127 0.013
R4815 a_6224_252.n58 a_6224_252.n57 0.008
R4816 a_6224_252.n125 a_6224_252.n124 0.008
R4817 VB.n6 VB.n5 1034.69
R4818 VB.n13 VB.n12 967.747
R4819 VB.n11 VB.t0 906.159
R4820 VB.n10 VB.n0 906.159
R4821 VB.n9 VB.n1 906.159
R4822 VB.n8 VB.n2 906.159
R4823 VB.n7 VB.n3 906.159
R4824 VB.n6 VB.n4 906.159
R4825 VB VB.n13 181.785
R4826 VB.n7 VB.n6 128.533
R4827 VB.n8 VB.n7 128.533
R4828 VB.n9 VB.n8 128.533
R4829 VB.n10 VB.n9 128.533
R4830 VB.n11 VB.n10 128.533
R4831 VB.n13 VB.n11 66.944
C0 VP VCT 6.94fF
C1 VP OUT 0.13fF
.ends

